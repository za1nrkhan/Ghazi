VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ghazi_top_dffram_csv
  CLASS BLOCK ;
  FOREIGN ghazi_top_dffram_csv ;
  ORIGIN 0.000 0.000 ;
  SIZE 2667.000 BY 3667.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3542.160 21.000 3542.760 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1691.200 2667.000 1691.800 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2001.530 3663.000 2001.810 3667.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.850 17.000 2251.130 21.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1831.280 21.000 1831.880 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 639.920 21.000 640.520 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.410 3663.000 105.690 3667.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 623.370 17.000 623.650 21.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.170 3663.000 1465.450 3667.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 53.760 2667.000 54.360 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 995.050 3663.000 995.330 3667.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1194.800 2667.000 1195.400 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 220.410 17.000 220.690 21.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1385.200 21.000 1385.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 572.770 17.000 573.050 21.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1950.930 3663.000 1951.210 3667.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 400.560 2667.000 401.160 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1037.040 21.000 1037.640 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 338.170 17.000 338.450 21.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1434.160 21.000 1434.760 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2956.000 2667.000 2956.600 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 673.970 17.000 674.250 21.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3145.040 21.000 3145.640 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2636.330 17.000 2636.610 21.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 978.490 3663.000 978.770 3667.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 367.920 21.000 368.520 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1112.810 3663.000 1113.090 3667.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 911.330 3663.000 911.610 3667.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1395.250 17.000 1395.530 21.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3029.440 2667.000 3030.040 ;
    END
  END io_in[36]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2555.370 3663.000 2555.650 3667.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2261.040 2667.000 2261.640 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.610 17.000 1126.890 21.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.930 17.000 456.210 21.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3600.640 2667.000 3601.240 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1414.570 3663.000 1414.850 3667.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.250 3663.000 38.530 3667.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 408.090 3663.000 408.370 3667.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2236.560 2667.000 2237.160 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3302.800 2667.000 3303.400 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1889.760 2667.000 1890.360 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 937.760 21.000 938.360 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 441.210 3663.000 441.490 3667.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 556.210 17.000 556.490 21.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 773.200 2667.000 773.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 765.040 21.000 765.640 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1839.440 2667.000 1840.040 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2183.690 17.000 2183.970 21.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 421.890 17.000 422.170 21.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.970 3663.000 559.250 3667.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3253.840 2667.000 3254.440 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.090 3663.000 1834.370 3667.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1814.960 2667.000 1815.560 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 317.600 21.000 318.200 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1483.120 21.000 1483.720 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2267.410 17.000 2267.690 21.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1814.770 17.000 1815.050 21.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3649.600 2667.000 3650.200 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2370.450 3663.000 2370.730 3667.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 104.080 2667.000 104.680 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1347.410 3663.000 1347.690 3667.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1409.680 21.000 1410.280 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1646.410 17.000 1646.690 21.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 21.690 3663.000 21.970 3667.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 3294.640 21.000 3295.240 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 472.490 17.000 472.770 21.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1608.240 21.000 1608.840 ;
    END
  END io_oeb[36]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 3467.360 21.000 3467.960 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2360.320 2667.000 2360.920 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 789.520 21.000 790.120 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2504.770 3663.000 2505.050 3667.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 659.250 3663.000 659.530 3667.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2639.090 3663.000 2639.370 3667.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1445.850 17.000 1446.130 21.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2102.730 3663.000 2103.010 3667.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 606.810 17.000 607.090 21.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 491.810 3663.000 492.090 3667.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.490 3663.000 357.770 3667.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 757.690 17.000 757.970 21.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2099.970 17.000 2100.250 21.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2200.250 17.000 2200.530 21.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2161.760 2667.000 2162.360 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3377.600 2667.000 3378.200 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2847.200 21.000 2847.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.970 17.000 53.250 21.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.050 17.000 305.330 21.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1532.330 3663.000 1532.610 3667.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 690.240 21.000 690.840 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1697.010 17.000 1697.290 21.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.730 17.000 355.010 21.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 723.650 17.000 723.930 21.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2452.330 17.000 2452.610 21.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2435.120 2667.000 2435.720 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2451.440 21.000 2452.040 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 590.250 17.000 590.530 21.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 508.370 3663.000 508.650 3667.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 656.490 17.000 656.770 21.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1632.720 21.000 1633.320 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3501.360 2667.000 3501.960 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1078.770 3663.000 1079.050 3667.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1020.720 2667.000 1021.320 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1598.570 3663.000 1598.850 3667.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 961.010 3663.000 961.290 3667.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 273.770 3663.000 274.050 3667.000 ;
    END
  END io_out[36]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1170.320 2667.000 1170.920 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1955.040 21.000 1955.640 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3451.040 2667.000 3451.640 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1649.170 3663.000 1649.450 3667.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1567.440 2667.000 1568.040 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1806.800 21.000 1807.400 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2169.890 3663.000 2170.170 3667.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 774.250 17.000 774.530 21.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1680.450 17.000 1680.730 21.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.890 3663.000 123.170 3667.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1462.410 17.000 1462.690 21.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 947.280 2667.000 947.880 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 475.360 2667.000 475.960 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 675.810 3663.000 676.090 3667.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2320.770 3663.000 2321.050 3667.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1699.770 3663.000 1700.050 3667.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2351.130 17.000 2351.410 21.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1359.360 21.000 1359.960 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1368.880 2667.000 1369.480 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.210 3663.000 2488.490 3667.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1160.800 21.000 1161.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2376.640 21.000 2377.240 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.530 17.000 69.810 21.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1136.320 21.000 1136.920 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2502.010 17.000 2502.290 21.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 29.280 2667.000 29.880 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 709.850 3663.000 710.130 3667.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1211.120 21.000 1211.720 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 489.050 17.000 489.330 21.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.810 3663.000 1918.090 3667.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1931.610 17.000 1931.890 21.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 203.850 17.000 204.130 21.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3319.120 21.000 3319.720 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 888.800 21.000 889.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2674.480 21.000 2675.080 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2550.720 21.000 2551.320 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1764.640 2667.000 1765.240 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 962.240 21.000 962.840 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 351.600 2667.000 352.200 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2931.520 2667.000 2932.120 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3442.880 21.000 3443.480 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2655.650 3663.000 2655.930 3667.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 790.810 17.000 791.090 21.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 741.130 17.000 741.410 21.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.770 3663.000 895.050 3667.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 119.040 21.000 119.640 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 237.890 17.000 238.170 21.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 457.770 3663.000 458.050 3667.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 128.560 2667.000 129.160 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2152.410 3663.000 2152.690 3667.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1145.840 2667.000 1146.440 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.650 17.000 1965.930 21.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.010 17.000 271.290 21.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3402.080 2667.000 3402.680 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2086.960 2667.000 2087.560 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2583.360 2667.000 2583.960 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 742.970 3663.000 743.250 3667.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2004.000 21.000 2004.600 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1120.000 2667.000 1120.600 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 626.130 3663.000 626.410 3667.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2252.880 21.000 2253.480 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 925.130 17.000 925.410 21.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3476.880 2667.000 3477.480 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1790.480 2667.000 1791.080 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 416.880 21.000 417.480 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2881.200 2667.000 2881.800 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1783.490 3663.000 1783.770 3667.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2650.000 21.000 2650.600 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3071.600 21.000 3072.200 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3104.240 2667.000 3104.840 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2732.960 2667.000 2733.560 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.450 17.000 254.730 21.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2723.440 21.000 2724.040 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1548.890 3663.000 1549.170 3667.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 293.120 21.000 293.720 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3021.280 21.000 3021.880 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1046.560 2667.000 1047.160 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1582.010 3663.000 1582.290 3667.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3268.800 21.000 3269.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 942.610 17.000 942.890 21.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2385.170 17.000 2385.450 21.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1817.530 3663.000 1817.810 3667.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.000 13.000 21.000 2420.040 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2806.400 2667.000 2807.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1235.600 21.000 1236.200 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.290 17.000 187.570 21.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2038.000 2667.000 2038.600 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1901.250 3663.000 1901.530 3667.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2521.330 3663.000 2521.610 3667.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3327.280 2667.000 3327.880 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3426.560 2667.000 3427.160 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2569.170 17.000 2569.450 21.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 276.800 2667.000 277.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2150.570 17.000 2150.850 21.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1111.840 21.000 1112.440 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1968.410 3663.000 1968.690 3667.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 574.640 2667.000 575.240 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2029.840 21.000 2030.440 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1884.690 3663.000 1884.970 3667.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 491.680 21.000 492.280 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1915.050 17.000 1915.330 21.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1715.680 2667.000 1716.280 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3096.080 21.000 3096.680 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2500.400 21.000 2501.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3550.320 2667.000 3550.920 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1565.450 3663.000 1565.730 3667.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2401.730 17.000 2402.010 21.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1557.920 21.000 1558.520 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3592.480 21.000 3593.080 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 324.370 3663.000 324.650 3667.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1160.650 17.000 1160.930 21.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1517.120 2667.000 1517.720 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 748.720 2667.000 749.320 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1087.360 21.000 1087.960 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2653.810 17.000 2654.090 21.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2335.840 2667.000 2336.440 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2368.610 17.000 2368.890 21.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 376.080 2667.000 376.680 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3353.120 2667.000 3353.720 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1095.330 3663.000 1095.610 3667.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 153.250 17.000 153.530 21.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1731.050 17.000 1731.330 21.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2873.040 21.000 2873.640 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1012.560 21.000 1013.160 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2334.570 17.000 2334.850 21.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 475.250 3663.000 475.530 3667.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 227.840 2667.000 228.440 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 844.170 3663.000 844.450 3667.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2236.130 3663.000 2236.410 3667.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 913.280 21.000 913.880 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1780.960 21.000 1781.560 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1193.770 17.000 1194.050 21.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 306.890 3663.000 307.170 3667.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1095.520 2667.000 1096.120 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2624.160 21.000 2624.760 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2065.930 17.000 2066.210 21.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2410.640 2667.000 2411.240 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1904.720 21.000 1905.320 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1428.370 17.000 1428.650 21.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 78.240 2667.000 78.840 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 525.680 2667.000 526.280 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.770 17.000 389.050 21.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 170.730 17.000 171.010 21.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1963.200 2667.000 1963.800 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 615.440 21.000 616.040 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.170 17.000 959.450 21.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2897.520 21.000 2898.120 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2798.240 21.000 2798.840 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2698.960 21.000 2699.560 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2437.610 3663.000 2437.890 3667.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1546.130 17.000 1546.410 21.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 3368.080 21.000 3368.680 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.210 17.000 1798.490 21.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2054.320 21.000 2054.920 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2303.290 3663.000 2303.570 3667.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3525.840 2667.000 3526.440 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2049.370 17.000 2049.650 21.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1541.600 2667.000 1542.200 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1938.720 2667.000 1939.320 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 392.400 21.000 393.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2277.360 21.000 2277.960 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 877.290 3663.000 877.570 3667.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.570 3663.000 172.850 3667.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 988.080 21.000 988.680 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 975.730 17.000 976.010 21.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1750.370 3663.000 1750.650 3667.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1071.040 2667.000 1071.640 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1478.970 17.000 1479.250 21.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2519.490 17.000 2519.770 21.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.570 17.000 287.850 21.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1431.130 3663.000 1431.410 3667.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1683.210 3663.000 1683.490 3667.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1177.210 17.000 1177.490 21.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 153.040 2667.000 153.640 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 542.410 3663.000 542.690 3667.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2167.130 17.000 2167.410 21.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2856.720 2667.000 2857.320 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1213.090 3663.000 1213.370 3667.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3154.560 2667.000 3155.160 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 575.530 3663.000 575.810 3667.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2178.080 21.000 2178.680 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1417.840 2667.000 1418.440 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1582.400 21.000 1583.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3278.320 2667.000 3278.920 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2285.520 2667.000 2286.120 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2202.560 21.000 2203.160 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1665.360 2667.000 1665.960 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 523.090 17.000 523.370 21.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1640.880 2667.000 1641.480 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2228.400 21.000 2229.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 169.360 21.000 169.960 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1934.370 3663.000 1934.650 3667.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 450.880 2667.000 451.480 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1219.280 2667.000 1219.880 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 872.480 2667.000 873.080 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1529.570 17.000 1529.850 21.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2682.640 2667.000 2683.240 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.850 3663.000 89.130 3667.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 3244.320 21.000 3244.920 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1210.330 17.000 1210.610 21.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2035.570 3663.000 2035.850 3667.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1850.650 3663.000 1850.930 3667.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2311.360 2667.000 2311.960 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 777.010 3663.000 777.290 3667.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 992.290 17.000 992.570 21.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1334.880 21.000 1335.480 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1229.650 3663.000 1229.930 3667.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2605.970 3663.000 2606.250 3667.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 206.610 3663.000 206.890 3667.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1513.010 17.000 1513.290 21.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 467.200 21.000 467.800 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1310.400 21.000 1311.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2972.320 21.000 2972.920 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1244.370 17.000 1244.650 21.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3079.760 2667.000 3080.360 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 714.720 21.000 715.320 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2186.450 3663.000 2186.730 3667.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1632.610 3663.000 1632.890 3667.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1468.160 2667.000 1468.760 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1361.210 17.000 1361.490 21.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 739.200 21.000 739.800 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2905.680 2667.000 2906.280 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 203.360 2667.000 203.960 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1498.290 3663.000 1498.570 3667.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2013.520 2667.000 2014.120 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 841.410 17.000 841.690 21.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1984.970 3663.000 1985.250 3667.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 218.320 21.000 218.920 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1982.210 17.000 1982.490 21.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1026.330 17.000 1026.610 21.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2032.810 17.000 2033.090 21.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2301.450 17.000 2301.730 21.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1162.490 3663.000 1162.770 3667.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 268.640 21.000 269.240 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2062.480 2667.000 2063.080 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2586.650 17.000 2586.930 21.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 599.120 2667.000 599.720 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 177.520 2667.000 178.120 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 726.410 3663.000 726.690 3667.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2538.810 3663.000 2539.090 3667.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1260.930 17.000 1261.210 21.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2418.290 17.000 2418.570 21.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.690 17.000 136.970 21.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1269.600 2667.000 1270.200 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 566.480 21.000 567.080 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1008.850 17.000 1009.130 21.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1865.370 17.000 1865.650 21.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2085.250 3663.000 2085.530 3667.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1732.000 21.000 1732.600 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2137.280 2667.000 2137.880 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1898.490 17.000 1898.770 21.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2575.200 21.000 2575.800 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2116.530 17.000 2116.810 21.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 94.560 21.000 95.160 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 3045.760 21.000 3046.360 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 3195.360 21.000 3195.960 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 516.160 21.000 516.760 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1914.240 2667.000 1914.840 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 793.570 3663.000 793.850 3667.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1863.920 2667.000 1864.520 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 252.320 2667.000 252.920 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.050 3663.000 190.330 3667.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.570 17.000 103.850 21.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2455.090 3663.000 2455.370 3667.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2353.890 3663.000 2354.170 3667.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3393.920 21.000 3394.520 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2524.880 21.000 2525.480 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2832.240 2667.000 2832.840 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1196.530 3663.000 1196.810 3667.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1059.450 17.000 1059.730 21.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1143.170 17.000 1143.450 21.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2212.080 2667.000 2212.680 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1740.160 2667.000 1740.760 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 120.130 17.000 120.410 21.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1311.530 17.000 1311.810 21.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2980.480 2667.000 2981.080 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1045.650 3663.000 1045.930 3667.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2484.080 2667.000 2484.680 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1062.210 3663.000 1062.490 3667.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1800.050 3663.000 1800.330 3667.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1998.770 17.000 1999.050 21.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1378.690 17.000 1378.970 21.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2996.800 21.000 2997.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 343.440 21.000 344.040 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 693.290 3663.000 693.570 3667.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1330.850 3663.000 1331.130 3667.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1294.080 2667.000 1294.680 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1186.640 21.000 1187.240 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 524.930 3663.000 525.210 3667.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1716.330 3663.000 1716.610 3667.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 540.640 21.000 541.240 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 649.440 2667.000 650.040 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1296.810 3663.000 1297.090 3667.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 327.120 2667.000 327.720 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3576.160 2667.000 3576.760 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 896.960 2667.000 897.560 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.450 17.000 438.730 21.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1285.920 21.000 1286.520 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2119.290 3663.000 2119.570 3667.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2468.890 17.000 2469.170 21.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1318.560 2667.000 1319.160 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1442.320 2667.000 1442.920 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2781.920 2667.000 2782.520 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.690 3663.000 1447.970 3667.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 590.960 21.000 591.560 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1930.560 21.000 1931.160 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.090 17.000 1328.370 21.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2112.800 2667.000 2113.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1398.010 3663.000 1398.290 3667.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 996.240 2667.000 996.840 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2475.920 21.000 2476.520 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2658.160 2667.000 2658.760 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1294.050 17.000 1294.330 21.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 857.970 17.000 858.250 21.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 550.160 2667.000 550.760 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1562.690 17.000 1562.970 21.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 822.160 2667.000 822.760 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1579.250 17.000 1579.530 21.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2083.410 17.000 2083.690 21.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.410 17.000 36.690 21.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2603.210 17.000 2603.490 21.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 426.400 2667.000 427.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.610 3663.000 390.890 3667.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.010 3663.000 156.290 3667.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3418.400 21.000 3419.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2352.160 21.000 2352.760 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1681.680 21.000 1682.280 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2707.120 2667.000 2707.720 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3179.040 2667.000 3179.640 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.730 3663.000 2287.010 3667.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2757.440 2667.000 2758.040 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3170.880 21.000 3171.480 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 698.400 2667.000 699.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2203.010 3663.000 2203.290 3667.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2558.880 2667.000 2559.480 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1492.640 2667.000 1493.240 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1280.250 3663.000 1280.530 3667.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1481.730 3663.000 1482.010 3667.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 810.130 3663.000 810.410 3667.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2135.850 3663.000 2136.130 3667.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1411.810 17.000 1412.090 21.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2384.800 2667.000 2385.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 290.330 3663.000 290.610 3667.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.930 3663.000 2572.210 3667.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.730 3663.000 240.010 3667.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1867.210 3663.000 1867.490 3667.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2749.280 21.000 2749.880 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1458.640 21.000 1459.240 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3055.280 2667.000 3055.880 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 340.930 3663.000 341.210 3667.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2773.760 21.000 2774.360 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1145.930 3663.000 1146.210 3667.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1629.850 17.000 1630.130 21.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1616.400 2667.000 1617.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2283.970 17.000 2284.250 21.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 707.090 17.000 707.370 21.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2337.330 3663.000 2337.610 3667.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2078.800 21.000 2079.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1880.240 21.000 1880.840 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3228.000 2667.000 3228.600 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 864.320 21.000 864.920 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2822.720 21.000 2823.320 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1766.930 3663.000 1767.210 3667.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2253.610 3663.000 2253.890 3667.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2946.480 21.000 2947.080 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1343.040 2667.000 1343.640 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 892.010 17.000 892.290 21.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1277.490 17.000 1277.770 21.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.650 3663.000 424.930 3667.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1263.690 3663.000 1263.970 3667.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2534.400 2667.000 2535.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 223.170 3663.000 223.450 3667.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2922.000 21.000 2922.600 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3493.200 21.000 3493.800 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 971.760 2667.000 972.360 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1514.850 3663.000 1515.130 3667.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 665.760 21.000 666.360 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1393.360 2667.000 1393.960 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3004.960 2667.000 3005.560 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2588.490 3663.000 2588.770 3667.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 722.880 2667.000 723.480 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2301.840 21.000 2302.440 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 624.960 2667.000 625.560 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 927.890 3663.000 928.170 3667.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 848.000 2667.000 848.600 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 639.930 17.000 640.210 21.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1533.440 21.000 1534.040 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2052.130 3663.000 2052.410 3667.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2552.610 17.000 2552.890 21.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1665.730 3663.000 1666.010 3667.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2485.450 17.000 2485.730 21.000 ;
    END
  END la_oen[9]
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 499.840 2667.000 500.440 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2129.120 21.000 2129.720 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2016.250 17.000 2016.530 21.000 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1110.050 17.000 1110.330 21.000 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3219.840 21.000 3220.440 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 944.450 3663.000 944.730 3667.000 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1657.200 21.000 1657.800 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3203.520 2667.000 3204.120 ;
    END
  END vssd2
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1713.570 17.000 1713.850 21.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 690.530 17.000 690.810 21.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1831.330 17.000 1831.610 21.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.730 3663.000 56.010 3667.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3343.600 21.000 3344.200 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1313.370 3663.000 1313.650 3667.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3566.640 21.000 3567.240 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2387.930 3663.000 2388.210 3667.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1732.890 3663.000 1733.170 3667.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1243.760 2667.000 1244.360 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1042.890 17.000 1043.170 21.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1508.960 21.000 1509.560 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1855.760 21.000 1856.360 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1260.080 21.000 1260.680 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.970 3663.000 1180.250 3667.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2471.650 3663.000 2471.930 3667.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1979.520 21.000 1980.120 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 244.160 21.000 244.760 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 673.920 2667.000 674.520 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2633.680 2667.000 2634.280 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1129.370 3663.000 1129.650 3667.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 609.570 3663.000 609.850 3667.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2607.840 2667.000 2608.440 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2133.090 17.000 2133.370 21.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 875.450 17.000 875.730 21.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 193.840 21.000 194.440 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1076.010 17.000 1076.290 21.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1247.130 3663.000 1247.410 3667.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2435.770 17.000 2436.050 21.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1591.920 2667.000 1592.520 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 442.720 21.000 443.320 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.930 17.000 1882.210 21.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1028.170 3663.000 1028.450 3667.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.730 17.000 1597.010 21.000 ;
    END
  END wbs_clk_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1847.890 17.000 1848.170 21.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 505.610 17.000 505.890 21.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 838.480 21.000 839.080 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2234.290 17.000 2234.570 21.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.450 3663.000 139.730 3667.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1344.650 17.000 1344.930 21.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 1756.480 21.000 1757.080 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2421.050 3663.000 2421.330 3667.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 144.880 21.000 145.480 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2404.490 3663.000 2404.770 3667.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3625.120 2667.000 3625.720 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2068.690 3663.000 2068.970 3667.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1093.490 17.000 1093.770 21.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.290 3663.000 72.570 3667.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2599.680 21.000 2600.280 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1363.970 3663.000 1364.250 3667.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2459.600 2667.000 2460.200 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2509.920 2667.000 2510.520 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3616.960 21.000 3617.560 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 908.570 17.000 908.850 21.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 797.680 2667.000 798.280 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 921.440 2667.000 922.040 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2318.010 17.000 2318.290 21.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.290 17.000 371.570 21.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 2186.240 2667.000 2186.840 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1747.610 17.000 1747.890 21.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1227.810 17.000 1228.090 21.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1764.170 17.000 1764.450 21.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2425.040 2533.640 2433.040 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2536.050 17.000 2536.330 21.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1380.530 3663.000 1380.810 3667.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 808.290 17.000 808.570 21.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 860.730 3663.000 861.010 3667.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2219.570 3663.000 2219.850 3667.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2103.280 21.000 2103.880 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1011.610 3663.000 1011.890 3667.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.770 17.000 2620.050 21.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1707.520 21.000 1708.120 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 301.280 2667.000 301.880 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.530 17.000 1495.810 21.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 1061.520 21.000 1062.120 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 3641.440 21.000 3642.040 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2622.530 3663.000 2622.810 3667.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1663.890 17.000 1664.170 21.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 321.610 17.000 321.890 21.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2270.170 3663.000 2270.450 3667.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 374.050 3663.000 374.330 3667.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 760.450 3663.000 760.730 3667.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 405.330 17.000 405.610 21.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 70.080 21.000 70.680 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 824.850 17.000 825.130 21.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1949.090 17.000 1949.370 21.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2216.810 17.000 2217.090 21.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2326.320 21.000 2326.920 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 592.090 3663.000 592.370 3667.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 45.600 21.000 46.200 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 2401.120 21.000 2401.720 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2663.000 3128.720 2667.000 3129.320 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 827.610 3663.000 827.890 3667.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.090 17.000 86.370 21.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 814.000 21.000 814.600 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 17.000 3517.680 21.000 3518.280 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 642.690 3663.000 642.970 3667.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2018.090 3663.000 2018.370 3667.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1616.050 3663.000 1616.330 3667.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_rst_ni
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 257.210 3663.000 257.490 3667.000 ;
    END
  END wbs_rst_ni
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1780.730 17.000 1781.010 21.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1613.290 17.000 1613.570 21.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 3120.560 21.000 3121.160 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.000 2153.600 21.000 2154.200 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2663.000 1989.040 2667.000 1989.640 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 539.650 17.000 539.930 21.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 17.000 32.610 2516.640 34.210 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 17.000 109.200 2516.640 110.800 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 17.000 16.915 2652.195 3643.355 ;
      LAYER met1 ;
        RECT 17.000 16.760 2652.730 3662.780 ;
      LAYER met2 ;
        RECT 0.000 3662.720 21.410 3663.000 ;
        RECT 22.250 3662.720 37.970 3663.000 ;
        RECT 38.810 3662.720 55.450 3663.000 ;
        RECT 56.290 3662.720 72.010 3663.000 ;
        RECT 72.850 3662.720 88.570 3663.000 ;
        RECT 89.410 3662.720 105.130 3663.000 ;
        RECT 105.970 3662.720 122.610 3663.000 ;
        RECT 123.450 3662.720 139.170 3663.000 ;
        RECT 140.010 3662.720 155.730 3663.000 ;
        RECT 156.570 3662.720 172.290 3663.000 ;
        RECT 173.130 3662.720 189.770 3663.000 ;
        RECT 190.610 3662.720 206.330 3663.000 ;
        RECT 207.170 3662.720 222.890 3663.000 ;
        RECT 223.730 3662.720 239.450 3663.000 ;
        RECT 240.290 3662.720 256.930 3663.000 ;
        RECT 257.770 3662.720 273.490 3663.000 ;
        RECT 274.330 3662.720 290.050 3663.000 ;
        RECT 290.890 3662.720 306.610 3663.000 ;
        RECT 307.450 3662.720 324.090 3663.000 ;
        RECT 324.930 3662.720 340.650 3663.000 ;
        RECT 341.490 3662.720 357.210 3663.000 ;
        RECT 358.050 3662.720 373.770 3663.000 ;
        RECT 374.610 3662.720 390.330 3663.000 ;
        RECT 391.170 3662.720 407.810 3663.000 ;
        RECT 408.650 3662.720 424.370 3663.000 ;
        RECT 425.210 3662.720 440.930 3663.000 ;
        RECT 441.770 3662.720 457.490 3663.000 ;
        RECT 458.330 3662.720 474.970 3663.000 ;
        RECT 475.810 3662.720 491.530 3663.000 ;
        RECT 492.370 3662.720 508.090 3663.000 ;
        RECT 508.930 3662.720 524.650 3663.000 ;
        RECT 525.490 3662.720 542.130 3663.000 ;
        RECT 542.970 3662.720 558.690 3663.000 ;
        RECT 559.530 3662.720 575.250 3663.000 ;
        RECT 576.090 3662.720 591.810 3663.000 ;
        RECT 592.650 3662.720 609.290 3663.000 ;
        RECT 610.130 3662.720 625.850 3663.000 ;
        RECT 626.690 3662.720 642.410 3663.000 ;
        RECT 643.250 3662.720 658.970 3663.000 ;
        RECT 659.810 3662.720 675.530 3663.000 ;
        RECT 676.370 3662.720 693.010 3663.000 ;
        RECT 693.850 3662.720 709.570 3663.000 ;
        RECT 710.410 3662.720 726.130 3663.000 ;
        RECT 726.970 3662.720 742.690 3663.000 ;
        RECT 743.530 3662.720 760.170 3663.000 ;
        RECT 761.010 3662.720 776.730 3663.000 ;
        RECT 777.570 3662.720 793.290 3663.000 ;
        RECT 794.130 3662.720 809.850 3663.000 ;
        RECT 810.690 3662.720 827.330 3663.000 ;
        RECT 828.170 3662.720 843.890 3663.000 ;
        RECT 844.730 3662.720 860.450 3663.000 ;
        RECT 861.290 3662.720 877.010 3663.000 ;
        RECT 877.850 3662.720 894.490 3663.000 ;
        RECT 895.330 3662.720 911.050 3663.000 ;
        RECT 911.890 3662.720 927.610 3663.000 ;
        RECT 928.450 3662.720 944.170 3663.000 ;
        RECT 945.010 3662.720 960.730 3663.000 ;
        RECT 961.570 3662.720 978.210 3663.000 ;
        RECT 979.050 3662.720 994.770 3663.000 ;
        RECT 995.610 3662.720 1011.330 3663.000 ;
        RECT 1012.170 3662.720 1027.890 3663.000 ;
        RECT 1028.730 3662.720 1045.370 3663.000 ;
        RECT 1046.210 3662.720 1061.930 3663.000 ;
        RECT 1062.770 3662.720 1078.490 3663.000 ;
        RECT 1079.330 3662.720 1095.050 3663.000 ;
        RECT 1095.890 3662.720 1112.530 3663.000 ;
        RECT 1113.370 3662.720 1129.090 3663.000 ;
        RECT 1129.930 3662.720 1145.650 3663.000 ;
        RECT 1146.490 3662.720 1162.210 3663.000 ;
        RECT 1163.050 3662.720 1179.690 3663.000 ;
        RECT 1180.530 3662.720 1196.250 3663.000 ;
        RECT 1197.090 3662.720 1212.810 3663.000 ;
        RECT 1213.650 3662.720 1229.370 3663.000 ;
        RECT 1230.210 3662.720 1246.850 3663.000 ;
        RECT 1247.690 3662.720 1263.410 3663.000 ;
        RECT 1264.250 3662.720 1279.970 3663.000 ;
        RECT 1280.810 3662.720 1296.530 3663.000 ;
        RECT 1297.370 3662.720 1313.090 3663.000 ;
        RECT 1313.930 3662.720 1330.570 3663.000 ;
        RECT 1331.410 3662.720 1347.130 3663.000 ;
        RECT 1347.970 3662.720 1363.690 3663.000 ;
        RECT 1364.530 3662.720 1380.250 3663.000 ;
        RECT 1381.090 3662.720 1397.730 3663.000 ;
        RECT 1398.570 3662.720 1414.290 3663.000 ;
        RECT 1415.130 3662.720 1430.850 3663.000 ;
        RECT 1431.690 3662.720 1447.410 3663.000 ;
        RECT 1448.250 3662.720 1464.890 3663.000 ;
        RECT 1465.730 3662.720 1481.450 3663.000 ;
        RECT 1482.290 3662.720 1498.010 3663.000 ;
        RECT 1498.850 3662.720 1514.570 3663.000 ;
        RECT 1515.410 3662.720 1532.050 3663.000 ;
        RECT 1532.890 3662.720 1548.610 3663.000 ;
        RECT 1549.450 3662.720 1565.170 3663.000 ;
        RECT 1566.010 3662.720 1581.730 3663.000 ;
        RECT 1582.570 3662.720 1598.290 3663.000 ;
        RECT 1599.130 3662.720 1615.770 3663.000 ;
        RECT 1616.610 3662.720 1632.330 3663.000 ;
        RECT 1633.170 3662.720 1648.890 3663.000 ;
        RECT 1649.730 3662.720 1665.450 3663.000 ;
        RECT 1666.290 3662.720 1682.930 3663.000 ;
        RECT 1683.770 3662.720 1699.490 3663.000 ;
        RECT 1700.330 3662.720 1716.050 3663.000 ;
        RECT 1716.890 3662.720 1732.610 3663.000 ;
        RECT 1733.450 3662.720 1750.090 3663.000 ;
        RECT 1750.930 3662.720 1766.650 3663.000 ;
        RECT 1767.490 3662.720 1783.210 3663.000 ;
        RECT 1784.050 3662.720 1799.770 3663.000 ;
        RECT 1800.610 3662.720 1817.250 3663.000 ;
        RECT 1818.090 3662.720 1833.810 3663.000 ;
        RECT 1834.650 3662.720 1850.370 3663.000 ;
        RECT 1851.210 3662.720 1866.930 3663.000 ;
        RECT 1867.770 3662.720 1884.410 3663.000 ;
        RECT 1885.250 3662.720 1900.970 3663.000 ;
        RECT 1901.810 3662.720 1917.530 3663.000 ;
        RECT 1918.370 3662.720 1934.090 3663.000 ;
        RECT 1934.930 3662.720 1950.650 3663.000 ;
        RECT 1951.490 3662.720 1968.130 3663.000 ;
        RECT 1968.970 3662.720 1984.690 3663.000 ;
        RECT 1985.530 3662.720 2001.250 3663.000 ;
        RECT 2002.090 3662.720 2017.810 3663.000 ;
        RECT 2018.650 3662.720 2035.290 3663.000 ;
        RECT 2036.130 3662.720 2051.850 3663.000 ;
        RECT 2052.690 3662.720 2068.410 3663.000 ;
        RECT 2069.250 3662.720 2084.970 3663.000 ;
        RECT 2085.810 3662.720 2102.450 3663.000 ;
        RECT 2103.290 3662.720 2119.010 3663.000 ;
        RECT 2119.850 3662.720 2135.570 3663.000 ;
        RECT 2136.410 3662.720 2152.130 3663.000 ;
        RECT 2152.970 3662.720 2169.610 3663.000 ;
        RECT 2170.450 3662.720 2186.170 3663.000 ;
        RECT 2187.010 3662.720 2202.730 3663.000 ;
        RECT 2203.570 3662.720 2219.290 3663.000 ;
        RECT 2220.130 3662.720 2235.850 3663.000 ;
        RECT 2236.690 3662.720 2253.330 3663.000 ;
        RECT 2254.170 3662.720 2269.890 3663.000 ;
        RECT 2270.730 3662.720 2286.450 3663.000 ;
        RECT 2287.290 3662.720 2303.010 3663.000 ;
        RECT 2303.850 3662.720 2320.490 3663.000 ;
        RECT 2321.330 3662.720 2337.050 3663.000 ;
        RECT 2337.890 3662.720 2353.610 3663.000 ;
        RECT 2354.450 3662.720 2370.170 3663.000 ;
        RECT 2371.010 3662.720 2387.650 3663.000 ;
        RECT 2388.490 3662.720 2404.210 3663.000 ;
        RECT 2405.050 3662.720 2420.770 3663.000 ;
        RECT 2421.610 3662.720 2437.330 3663.000 ;
        RECT 2438.170 3662.720 2454.810 3663.000 ;
        RECT 2455.650 3662.720 2471.370 3663.000 ;
        RECT 2472.210 3662.720 2487.930 3663.000 ;
        RECT 2488.770 3662.720 2504.490 3663.000 ;
        RECT 2505.330 3662.720 2521.050 3663.000 ;
        RECT 2521.890 3662.720 2538.530 3663.000 ;
        RECT 2539.370 3662.720 2555.090 3663.000 ;
        RECT 2555.930 3662.720 2571.650 3663.000 ;
        RECT 2572.490 3662.720 2588.210 3663.000 ;
        RECT 2589.050 3662.720 2605.690 3663.000 ;
        RECT 2606.530 3662.720 2622.250 3663.000 ;
        RECT 2623.090 3662.720 2638.810 3663.000 ;
        RECT 2639.650 3662.720 2655.370 3663.000 ;
        RECT 0.000 2420.320 2655.930 3662.720 ;
        RECT 0.000 12.720 12.720 2420.320 ;
        RECT 21.280 21.280 2655.930 2420.320 ;
        RECT 21.280 16.720 36.130 21.280 ;
        RECT 36.970 16.720 52.690 21.280 ;
        RECT 53.530 16.720 69.250 21.280 ;
        RECT 70.090 16.720 85.810 21.280 ;
        RECT 86.650 16.720 103.290 21.280 ;
        RECT 104.130 16.720 119.850 21.280 ;
        RECT 120.690 16.720 136.410 21.280 ;
        RECT 137.250 16.720 152.970 21.280 ;
        RECT 153.810 16.720 170.450 21.280 ;
        RECT 171.290 16.720 187.010 21.280 ;
        RECT 187.850 16.720 203.570 21.280 ;
        RECT 204.410 16.720 220.130 21.280 ;
        RECT 220.970 16.720 237.610 21.280 ;
        RECT 238.450 16.720 254.170 21.280 ;
        RECT 255.010 16.720 270.730 21.280 ;
        RECT 271.570 16.720 287.290 21.280 ;
        RECT 288.130 16.720 304.770 21.280 ;
        RECT 305.610 16.720 321.330 21.280 ;
        RECT 322.170 16.720 337.890 21.280 ;
        RECT 338.730 16.720 354.450 21.280 ;
        RECT 355.290 16.720 371.010 21.280 ;
        RECT 371.850 16.720 388.490 21.280 ;
        RECT 389.330 16.720 405.050 21.280 ;
        RECT 405.890 16.720 421.610 21.280 ;
        RECT 422.450 16.720 438.170 21.280 ;
        RECT 439.010 16.720 455.650 21.280 ;
        RECT 456.490 16.720 472.210 21.280 ;
        RECT 473.050 16.720 488.770 21.280 ;
        RECT 489.610 16.720 505.330 21.280 ;
        RECT 506.170 16.720 522.810 21.280 ;
        RECT 523.650 16.720 539.370 21.280 ;
        RECT 540.210 16.720 555.930 21.280 ;
        RECT 556.770 16.720 572.490 21.280 ;
        RECT 573.330 16.720 589.970 21.280 ;
        RECT 590.810 16.720 606.530 21.280 ;
        RECT 607.370 16.720 623.090 21.280 ;
        RECT 623.930 16.720 639.650 21.280 ;
        RECT 640.490 16.720 656.210 21.280 ;
        RECT 657.050 16.720 673.690 21.280 ;
        RECT 674.530 16.720 690.250 21.280 ;
        RECT 691.090 16.720 706.810 21.280 ;
        RECT 707.650 16.720 723.370 21.280 ;
        RECT 724.210 16.720 740.850 21.280 ;
        RECT 741.690 16.720 757.410 21.280 ;
        RECT 758.250 16.720 773.970 21.280 ;
        RECT 774.810 16.720 790.530 21.280 ;
        RECT 791.370 16.720 808.010 21.280 ;
        RECT 808.850 16.720 824.570 21.280 ;
        RECT 825.410 16.720 841.130 21.280 ;
        RECT 841.970 16.720 857.690 21.280 ;
        RECT 858.530 16.720 875.170 21.280 ;
        RECT 876.010 16.720 891.730 21.280 ;
        RECT 892.570 16.720 908.290 21.280 ;
        RECT 909.130 16.720 924.850 21.280 ;
        RECT 925.690 16.720 942.330 21.280 ;
        RECT 943.170 16.720 958.890 21.280 ;
        RECT 959.730 16.720 975.450 21.280 ;
        RECT 976.290 16.720 992.010 21.280 ;
        RECT 992.850 16.720 1008.570 21.280 ;
        RECT 1009.410 16.720 1026.050 21.280 ;
        RECT 1026.890 16.720 1042.610 21.280 ;
        RECT 1043.450 16.720 1059.170 21.280 ;
        RECT 1060.010 16.720 1075.730 21.280 ;
        RECT 1076.570 16.720 1093.210 21.280 ;
        RECT 1094.050 16.720 1109.770 21.280 ;
        RECT 1110.610 16.720 1126.330 21.280 ;
        RECT 1127.170 16.720 1142.890 21.280 ;
        RECT 1143.730 16.720 1160.370 21.280 ;
        RECT 1161.210 16.720 1176.930 21.280 ;
        RECT 1177.770 16.720 1193.490 21.280 ;
        RECT 1194.330 16.720 1210.050 21.280 ;
        RECT 1210.890 16.720 1227.530 21.280 ;
        RECT 1228.370 16.720 1244.090 21.280 ;
        RECT 1244.930 16.720 1260.650 21.280 ;
        RECT 1261.490 16.720 1277.210 21.280 ;
        RECT 1278.050 16.720 1293.770 21.280 ;
        RECT 1294.610 16.720 1311.250 21.280 ;
        RECT 1312.090 16.720 1327.810 21.280 ;
        RECT 1328.650 16.720 1344.370 21.280 ;
        RECT 1345.210 16.720 1360.930 21.280 ;
        RECT 1361.770 16.720 1378.410 21.280 ;
        RECT 1379.250 16.720 1394.970 21.280 ;
        RECT 1395.810 16.720 1411.530 21.280 ;
        RECT 1412.370 16.720 1428.090 21.280 ;
        RECT 1428.930 16.720 1445.570 21.280 ;
        RECT 1446.410 16.720 1462.130 21.280 ;
        RECT 1462.970 16.720 1478.690 21.280 ;
        RECT 1479.530 16.720 1495.250 21.280 ;
        RECT 1496.090 16.720 1512.730 21.280 ;
        RECT 1513.570 16.720 1529.290 21.280 ;
        RECT 1530.130 16.720 1545.850 21.280 ;
        RECT 1546.690 16.720 1562.410 21.280 ;
        RECT 1563.250 16.720 1578.970 21.280 ;
        RECT 1579.810 16.720 1596.450 21.280 ;
        RECT 1597.290 16.720 1613.010 21.280 ;
        RECT 1613.850 16.720 1629.570 21.280 ;
        RECT 1630.410 16.720 1646.130 21.280 ;
        RECT 1646.970 16.720 1663.610 21.280 ;
        RECT 1664.450 16.720 1680.170 21.280 ;
        RECT 1681.010 16.720 1696.730 21.280 ;
        RECT 1697.570 16.720 1713.290 21.280 ;
        RECT 1714.130 16.720 1730.770 21.280 ;
        RECT 1731.610 16.720 1747.330 21.280 ;
        RECT 1748.170 16.720 1763.890 21.280 ;
        RECT 1764.730 16.720 1780.450 21.280 ;
        RECT 1781.290 16.720 1797.930 21.280 ;
        RECT 1798.770 16.720 1814.490 21.280 ;
        RECT 1815.330 16.720 1831.050 21.280 ;
        RECT 1831.890 16.720 1847.610 21.280 ;
        RECT 1848.450 16.720 1865.090 21.280 ;
        RECT 1865.930 16.720 1881.650 21.280 ;
        RECT 1882.490 16.720 1898.210 21.280 ;
        RECT 1899.050 16.720 1914.770 21.280 ;
        RECT 1915.610 16.720 1931.330 21.280 ;
        RECT 1932.170 16.720 1948.810 21.280 ;
        RECT 1949.650 16.720 1965.370 21.280 ;
        RECT 1966.210 16.720 1981.930 21.280 ;
        RECT 1982.770 16.720 1998.490 21.280 ;
        RECT 1999.330 16.720 2015.970 21.280 ;
        RECT 2016.810 16.720 2032.530 21.280 ;
        RECT 2033.370 16.720 2049.090 21.280 ;
        RECT 2049.930 16.720 2065.650 21.280 ;
        RECT 2066.490 16.720 2083.130 21.280 ;
        RECT 2083.970 16.720 2099.690 21.280 ;
        RECT 2100.530 16.720 2116.250 21.280 ;
        RECT 2117.090 16.720 2132.810 21.280 ;
        RECT 2133.650 16.720 2150.290 21.280 ;
        RECT 2151.130 16.720 2166.850 21.280 ;
        RECT 2167.690 16.720 2183.410 21.280 ;
        RECT 2184.250 16.720 2199.970 21.280 ;
        RECT 2200.810 16.720 2216.530 21.280 ;
        RECT 2217.370 16.720 2234.010 21.280 ;
        RECT 2234.850 16.720 2250.570 21.280 ;
        RECT 2251.410 16.720 2267.130 21.280 ;
        RECT 2267.970 16.720 2283.690 21.280 ;
        RECT 2284.530 16.720 2301.170 21.280 ;
        RECT 2302.010 16.720 2317.730 21.280 ;
        RECT 2318.570 16.720 2334.290 21.280 ;
        RECT 2335.130 16.720 2350.850 21.280 ;
        RECT 2351.690 16.720 2368.330 21.280 ;
        RECT 2369.170 16.720 2384.890 21.280 ;
        RECT 2385.730 16.720 2401.450 21.280 ;
        RECT 2402.290 16.720 2418.010 21.280 ;
        RECT 2418.850 16.720 2435.490 21.280 ;
        RECT 2436.330 16.720 2452.050 21.280 ;
        RECT 2452.890 16.720 2468.610 21.280 ;
        RECT 2469.450 16.720 2485.170 21.280 ;
        RECT 2486.010 16.720 2501.730 21.280 ;
        RECT 2502.570 16.720 2519.210 21.280 ;
        RECT 2520.050 16.720 2535.770 21.280 ;
        RECT 2536.610 16.720 2552.330 21.280 ;
        RECT 2553.170 16.720 2568.890 21.280 ;
        RECT 2569.730 16.720 2586.370 21.280 ;
        RECT 2587.210 16.720 2602.930 21.280 ;
        RECT 2603.770 16.720 2619.490 21.280 ;
        RECT 2620.330 16.720 2636.050 21.280 ;
        RECT 2636.890 16.720 2653.530 21.280 ;
        RECT 2654.370 16.720 2655.930 21.280 ;
        RECT 21.280 12.720 2655.930 16.720 ;
        RECT 0.000 0.000 2655.930 12.720 ;
      LAYER met3 ;
        RECT 0.000 3649.200 2662.600 3650.065 ;
        RECT 0.000 3642.440 2663.000 3649.200 ;
        RECT 0.000 3641.040 16.600 3642.440 ;
        RECT 21.400 3641.040 2663.000 3642.440 ;
        RECT 0.000 3626.120 2663.000 3641.040 ;
        RECT 0.000 3624.720 2662.600 3626.120 ;
        RECT 0.000 3617.960 2663.000 3624.720 ;
        RECT 0.000 3616.560 16.600 3617.960 ;
        RECT 21.400 3616.560 2663.000 3617.960 ;
        RECT 0.000 3601.640 2663.000 3616.560 ;
        RECT 0.000 3600.240 2662.600 3601.640 ;
        RECT 0.000 3593.480 2663.000 3600.240 ;
        RECT 0.000 3592.080 16.600 3593.480 ;
        RECT 21.400 3592.080 2663.000 3593.480 ;
        RECT 0.000 3577.160 2663.000 3592.080 ;
        RECT 0.000 3575.760 2662.600 3577.160 ;
        RECT 0.000 3567.640 2663.000 3575.760 ;
        RECT 0.000 3566.240 16.600 3567.640 ;
        RECT 21.400 3566.240 2663.000 3567.640 ;
        RECT 0.000 3551.320 2663.000 3566.240 ;
        RECT 0.000 3549.920 2662.600 3551.320 ;
        RECT 0.000 3543.160 2663.000 3549.920 ;
        RECT 0.000 3541.760 16.600 3543.160 ;
        RECT 21.400 3541.760 2663.000 3543.160 ;
        RECT 0.000 3526.840 2663.000 3541.760 ;
        RECT 0.000 3525.440 2662.600 3526.840 ;
        RECT 0.000 3518.680 2663.000 3525.440 ;
        RECT 0.000 3517.280 16.600 3518.680 ;
        RECT 21.400 3517.280 2663.000 3518.680 ;
        RECT 0.000 3502.360 2663.000 3517.280 ;
        RECT 0.000 3500.960 2662.600 3502.360 ;
        RECT 0.000 3494.200 2663.000 3500.960 ;
        RECT 0.000 3492.800 16.600 3494.200 ;
        RECT 21.400 3492.800 2663.000 3494.200 ;
        RECT 0.000 3477.880 2663.000 3492.800 ;
        RECT 0.000 3476.480 2662.600 3477.880 ;
        RECT 0.000 3468.360 2663.000 3476.480 ;
        RECT 0.000 3466.960 16.600 3468.360 ;
        RECT 21.400 3466.960 2663.000 3468.360 ;
        RECT 0.000 3452.040 2663.000 3466.960 ;
        RECT 0.000 3450.640 2662.600 3452.040 ;
        RECT 0.000 3443.880 2663.000 3450.640 ;
        RECT 0.000 3442.480 16.600 3443.880 ;
        RECT 21.400 3442.480 2663.000 3443.880 ;
        RECT 0.000 3427.560 2663.000 3442.480 ;
        RECT 0.000 3426.160 2662.600 3427.560 ;
        RECT 0.000 3419.400 2663.000 3426.160 ;
        RECT 0.000 3418.000 16.600 3419.400 ;
        RECT 21.400 3418.000 2663.000 3419.400 ;
        RECT 0.000 3403.080 2663.000 3418.000 ;
        RECT 0.000 3401.680 2662.600 3403.080 ;
        RECT 0.000 3394.920 2663.000 3401.680 ;
        RECT 0.000 3393.520 16.600 3394.920 ;
        RECT 21.400 3393.520 2663.000 3394.920 ;
        RECT 0.000 3378.600 2663.000 3393.520 ;
        RECT 0.000 3377.200 2662.600 3378.600 ;
        RECT 0.000 3369.080 2663.000 3377.200 ;
        RECT 0.000 3367.680 16.600 3369.080 ;
        RECT 21.400 3367.680 2663.000 3369.080 ;
        RECT 0.000 3354.120 2663.000 3367.680 ;
        RECT 0.000 3352.720 2662.600 3354.120 ;
        RECT 0.000 3344.600 2663.000 3352.720 ;
        RECT 0.000 3343.200 16.600 3344.600 ;
        RECT 21.400 3343.200 2663.000 3344.600 ;
        RECT 0.000 3328.280 2663.000 3343.200 ;
        RECT 0.000 3326.880 2662.600 3328.280 ;
        RECT 0.000 3320.120 2663.000 3326.880 ;
        RECT 0.000 3318.720 16.600 3320.120 ;
        RECT 21.400 3318.720 2663.000 3320.120 ;
        RECT 0.000 3303.800 2663.000 3318.720 ;
        RECT 0.000 3302.400 2662.600 3303.800 ;
        RECT 0.000 3295.640 2663.000 3302.400 ;
        RECT 0.000 3294.240 16.600 3295.640 ;
        RECT 21.400 3294.240 2663.000 3295.640 ;
        RECT 0.000 3279.320 2663.000 3294.240 ;
        RECT 0.000 3277.920 2662.600 3279.320 ;
        RECT 0.000 3269.800 2663.000 3277.920 ;
        RECT 0.000 3268.400 16.600 3269.800 ;
        RECT 21.400 3268.400 2663.000 3269.800 ;
        RECT 0.000 3254.840 2663.000 3268.400 ;
        RECT 0.000 3253.440 2662.600 3254.840 ;
        RECT 0.000 3245.320 2663.000 3253.440 ;
        RECT 0.000 3243.920 16.600 3245.320 ;
        RECT 21.400 3243.920 2663.000 3245.320 ;
        RECT 0.000 3229.000 2663.000 3243.920 ;
        RECT 0.000 3227.600 2662.600 3229.000 ;
        RECT 0.000 3220.840 2663.000 3227.600 ;
        RECT 0.000 3219.440 16.600 3220.840 ;
        RECT 21.400 3219.440 2663.000 3220.840 ;
        RECT 0.000 3204.520 2663.000 3219.440 ;
        RECT 0.000 3203.120 2662.600 3204.520 ;
        RECT 0.000 3196.360 2663.000 3203.120 ;
        RECT 0.000 3194.960 16.600 3196.360 ;
        RECT 21.400 3194.960 2663.000 3196.360 ;
        RECT 0.000 3180.040 2663.000 3194.960 ;
        RECT 0.000 3178.640 2662.600 3180.040 ;
        RECT 0.000 3171.880 2663.000 3178.640 ;
        RECT 0.000 3170.480 16.600 3171.880 ;
        RECT 21.400 3170.480 2663.000 3171.880 ;
        RECT 0.000 3155.560 2663.000 3170.480 ;
        RECT 0.000 3154.160 2662.600 3155.560 ;
        RECT 0.000 3146.040 2663.000 3154.160 ;
        RECT 0.000 3144.640 16.600 3146.040 ;
        RECT 21.400 3144.640 2663.000 3146.040 ;
        RECT 0.000 3129.720 2663.000 3144.640 ;
        RECT 0.000 3128.320 2662.600 3129.720 ;
        RECT 0.000 3121.560 2663.000 3128.320 ;
        RECT 0.000 3120.160 16.600 3121.560 ;
        RECT 21.400 3120.160 2663.000 3121.560 ;
        RECT 0.000 3105.240 2663.000 3120.160 ;
        RECT 0.000 3103.840 2662.600 3105.240 ;
        RECT 0.000 3097.080 2663.000 3103.840 ;
        RECT 0.000 3095.680 16.600 3097.080 ;
        RECT 21.400 3095.680 2663.000 3097.080 ;
        RECT 0.000 3080.760 2663.000 3095.680 ;
        RECT 0.000 3079.360 2662.600 3080.760 ;
        RECT 0.000 3072.600 2663.000 3079.360 ;
        RECT 0.000 3071.200 16.600 3072.600 ;
        RECT 21.400 3071.200 2663.000 3072.600 ;
        RECT 0.000 3056.280 2663.000 3071.200 ;
        RECT 0.000 3054.880 2662.600 3056.280 ;
        RECT 0.000 3046.760 2663.000 3054.880 ;
        RECT 0.000 3045.360 16.600 3046.760 ;
        RECT 21.400 3045.360 2663.000 3046.760 ;
        RECT 0.000 3030.440 2663.000 3045.360 ;
        RECT 0.000 3029.040 2662.600 3030.440 ;
        RECT 0.000 3022.280 2663.000 3029.040 ;
        RECT 0.000 3020.880 16.600 3022.280 ;
        RECT 21.400 3020.880 2663.000 3022.280 ;
        RECT 0.000 3005.960 2663.000 3020.880 ;
        RECT 0.000 3004.560 2662.600 3005.960 ;
        RECT 0.000 2997.800 2663.000 3004.560 ;
        RECT 0.000 2996.400 16.600 2997.800 ;
        RECT 21.400 2996.400 2663.000 2997.800 ;
        RECT 0.000 2981.480 2663.000 2996.400 ;
        RECT 0.000 2980.080 2662.600 2981.480 ;
        RECT 0.000 2973.320 2663.000 2980.080 ;
        RECT 0.000 2971.920 16.600 2973.320 ;
        RECT 21.400 2971.920 2663.000 2973.320 ;
        RECT 0.000 2957.000 2663.000 2971.920 ;
        RECT 0.000 2955.600 2662.600 2957.000 ;
        RECT 0.000 2947.480 2663.000 2955.600 ;
        RECT 0.000 2946.080 16.600 2947.480 ;
        RECT 21.400 2946.080 2663.000 2947.480 ;
        RECT 0.000 2932.520 2663.000 2946.080 ;
        RECT 0.000 2931.120 2662.600 2932.520 ;
        RECT 0.000 2923.000 2663.000 2931.120 ;
        RECT 0.000 2921.600 16.600 2923.000 ;
        RECT 21.400 2921.600 2663.000 2923.000 ;
        RECT 0.000 2906.680 2663.000 2921.600 ;
        RECT 0.000 2905.280 2662.600 2906.680 ;
        RECT 0.000 2898.520 2663.000 2905.280 ;
        RECT 0.000 2897.120 16.600 2898.520 ;
        RECT 21.400 2897.120 2663.000 2898.520 ;
        RECT 0.000 2882.200 2663.000 2897.120 ;
        RECT 0.000 2880.800 2662.600 2882.200 ;
        RECT 0.000 2874.040 2663.000 2880.800 ;
        RECT 0.000 2872.640 16.600 2874.040 ;
        RECT 21.400 2872.640 2663.000 2874.040 ;
        RECT 0.000 2857.720 2663.000 2872.640 ;
        RECT 0.000 2856.320 2662.600 2857.720 ;
        RECT 0.000 2848.200 2663.000 2856.320 ;
        RECT 0.000 2846.800 16.600 2848.200 ;
        RECT 21.400 2846.800 2663.000 2848.200 ;
        RECT 0.000 2833.240 2663.000 2846.800 ;
        RECT 0.000 2831.840 2662.600 2833.240 ;
        RECT 0.000 2823.720 2663.000 2831.840 ;
        RECT 0.000 2822.320 16.600 2823.720 ;
        RECT 21.400 2822.320 2663.000 2823.720 ;
        RECT 0.000 2807.400 2663.000 2822.320 ;
        RECT 0.000 2806.000 2662.600 2807.400 ;
        RECT 0.000 2799.240 2663.000 2806.000 ;
        RECT 0.000 2797.840 16.600 2799.240 ;
        RECT 21.400 2797.840 2663.000 2799.240 ;
        RECT 0.000 2782.920 2663.000 2797.840 ;
        RECT 0.000 2781.520 2662.600 2782.920 ;
        RECT 0.000 2774.760 2663.000 2781.520 ;
        RECT 0.000 2773.360 16.600 2774.760 ;
        RECT 21.400 2773.360 2663.000 2774.760 ;
        RECT 0.000 2758.440 2663.000 2773.360 ;
        RECT 0.000 2757.040 2662.600 2758.440 ;
        RECT 0.000 2750.280 2663.000 2757.040 ;
        RECT 0.000 2748.880 16.600 2750.280 ;
        RECT 21.400 2748.880 2663.000 2750.280 ;
        RECT 0.000 2733.960 2663.000 2748.880 ;
        RECT 0.000 2732.560 2662.600 2733.960 ;
        RECT 0.000 2724.440 2663.000 2732.560 ;
        RECT 0.000 2723.040 16.600 2724.440 ;
        RECT 21.400 2723.040 2663.000 2724.440 ;
        RECT 0.000 2708.120 2663.000 2723.040 ;
        RECT 0.000 2706.720 2662.600 2708.120 ;
        RECT 0.000 2699.960 2663.000 2706.720 ;
        RECT 0.000 2698.560 16.600 2699.960 ;
        RECT 21.400 2698.560 2663.000 2699.960 ;
        RECT 0.000 2683.640 2663.000 2698.560 ;
        RECT 0.000 2682.240 2662.600 2683.640 ;
        RECT 0.000 2675.480 2663.000 2682.240 ;
        RECT 0.000 2674.080 16.600 2675.480 ;
        RECT 21.400 2674.080 2663.000 2675.480 ;
        RECT 0.000 2659.160 2663.000 2674.080 ;
        RECT 0.000 2657.760 2662.600 2659.160 ;
        RECT 0.000 2651.000 2663.000 2657.760 ;
        RECT 0.000 2649.600 16.600 2651.000 ;
        RECT 21.400 2649.600 2663.000 2651.000 ;
        RECT 0.000 2634.680 2663.000 2649.600 ;
        RECT 0.000 2633.280 2662.600 2634.680 ;
        RECT 0.000 2625.160 2663.000 2633.280 ;
        RECT 0.000 2623.760 16.600 2625.160 ;
        RECT 21.400 2623.760 2663.000 2625.160 ;
        RECT 0.000 2608.840 2663.000 2623.760 ;
        RECT 0.000 2607.440 2662.600 2608.840 ;
        RECT 0.000 2600.680 2663.000 2607.440 ;
        RECT 0.000 2599.280 16.600 2600.680 ;
        RECT 21.400 2599.280 2663.000 2600.680 ;
        RECT 0.000 2584.360 2663.000 2599.280 ;
        RECT 0.000 2582.960 2662.600 2584.360 ;
        RECT 0.000 2576.200 2663.000 2582.960 ;
        RECT 0.000 2574.800 16.600 2576.200 ;
        RECT 21.400 2574.800 2663.000 2576.200 ;
        RECT 0.000 2559.880 2663.000 2574.800 ;
        RECT 0.000 2558.480 2662.600 2559.880 ;
        RECT 0.000 2551.720 2663.000 2558.480 ;
        RECT 0.000 2550.320 16.600 2551.720 ;
        RECT 21.400 2550.320 2663.000 2551.720 ;
        RECT 0.000 2535.400 2663.000 2550.320 ;
        RECT 0.000 2534.000 2662.600 2535.400 ;
        RECT 0.000 2525.880 2663.000 2534.000 ;
        RECT 0.000 2524.480 16.600 2525.880 ;
        RECT 21.400 2524.480 2663.000 2525.880 ;
        RECT 0.000 2510.920 2663.000 2524.480 ;
        RECT 0.000 2509.520 2662.600 2510.920 ;
        RECT 0.000 2501.400 2663.000 2509.520 ;
        RECT 0.000 2500.000 16.600 2501.400 ;
        RECT 21.400 2500.000 2663.000 2501.400 ;
        RECT 0.000 2485.080 2663.000 2500.000 ;
        RECT 0.000 2483.680 2662.600 2485.080 ;
        RECT 0.000 2476.920 2663.000 2483.680 ;
        RECT 0.000 2475.520 16.600 2476.920 ;
        RECT 21.400 2475.520 2663.000 2476.920 ;
        RECT 0.000 2460.600 2663.000 2475.520 ;
        RECT 0.000 2459.200 2662.600 2460.600 ;
        RECT 0.000 2452.440 2663.000 2459.200 ;
        RECT 0.000 2451.040 16.600 2452.440 ;
        RECT 21.400 2451.040 2663.000 2452.440 ;
        RECT 0.000 2436.120 2663.000 2451.040 ;
        RECT 0.000 2434.720 2662.600 2436.120 ;
        RECT 0.000 2433.440 2663.000 2434.720 ;
        RECT 2534.040 2424.640 2663.000 2433.440 ;
        RECT 0.000 2411.640 2663.000 2424.640 ;
        RECT 0.000 2410.240 2662.600 2411.640 ;
        RECT 0.000 2402.120 2663.000 2410.240 ;
        RECT 0.000 2400.720 16.600 2402.120 ;
        RECT 21.400 2400.720 2663.000 2402.120 ;
        RECT 0.000 2385.800 2663.000 2400.720 ;
        RECT 0.000 2384.400 2662.600 2385.800 ;
        RECT 0.000 2377.640 2663.000 2384.400 ;
        RECT 0.000 2376.240 16.600 2377.640 ;
        RECT 21.400 2376.240 2663.000 2377.640 ;
        RECT 0.000 2361.320 2663.000 2376.240 ;
        RECT 0.000 2359.920 2662.600 2361.320 ;
        RECT 0.000 2353.160 2663.000 2359.920 ;
        RECT 0.000 2351.760 16.600 2353.160 ;
        RECT 21.400 2351.760 2663.000 2353.160 ;
        RECT 0.000 2336.840 2663.000 2351.760 ;
        RECT 0.000 2335.440 2662.600 2336.840 ;
        RECT 0.000 2327.320 2663.000 2335.440 ;
        RECT 0.000 2325.920 16.600 2327.320 ;
        RECT 21.400 2325.920 2663.000 2327.320 ;
        RECT 0.000 2312.360 2663.000 2325.920 ;
        RECT 0.000 2310.960 2662.600 2312.360 ;
        RECT 0.000 2302.840 2663.000 2310.960 ;
        RECT 0.000 2301.440 16.600 2302.840 ;
        RECT 21.400 2301.440 2663.000 2302.840 ;
        RECT 0.000 2286.520 2663.000 2301.440 ;
        RECT 0.000 2285.120 2662.600 2286.520 ;
        RECT 0.000 2278.360 2663.000 2285.120 ;
        RECT 0.000 2276.960 16.600 2278.360 ;
        RECT 21.400 2276.960 2663.000 2278.360 ;
        RECT 0.000 2262.040 2663.000 2276.960 ;
        RECT 0.000 2260.640 2662.600 2262.040 ;
        RECT 0.000 2253.880 2663.000 2260.640 ;
        RECT 0.000 2252.480 16.600 2253.880 ;
        RECT 21.400 2252.480 2663.000 2253.880 ;
        RECT 0.000 2237.560 2663.000 2252.480 ;
        RECT 0.000 2236.160 2662.600 2237.560 ;
        RECT 0.000 2229.400 2663.000 2236.160 ;
        RECT 0.000 2228.000 16.600 2229.400 ;
        RECT 21.400 2228.000 2663.000 2229.400 ;
        RECT 0.000 2213.080 2663.000 2228.000 ;
        RECT 0.000 2211.680 2662.600 2213.080 ;
        RECT 0.000 2203.560 2663.000 2211.680 ;
        RECT 0.000 2202.160 16.600 2203.560 ;
        RECT 21.400 2202.160 2663.000 2203.560 ;
        RECT 0.000 2187.240 2663.000 2202.160 ;
        RECT 0.000 2185.840 2662.600 2187.240 ;
        RECT 0.000 2179.080 2663.000 2185.840 ;
        RECT 0.000 2177.680 16.600 2179.080 ;
        RECT 21.400 2177.680 2663.000 2179.080 ;
        RECT 0.000 2162.760 2663.000 2177.680 ;
        RECT 0.000 2161.360 2662.600 2162.760 ;
        RECT 0.000 2154.600 2663.000 2161.360 ;
        RECT 0.000 2153.200 16.600 2154.600 ;
        RECT 21.400 2153.200 2663.000 2154.600 ;
        RECT 0.000 2138.280 2663.000 2153.200 ;
        RECT 0.000 2136.880 2662.600 2138.280 ;
        RECT 0.000 2130.120 2663.000 2136.880 ;
        RECT 0.000 2128.720 16.600 2130.120 ;
        RECT 21.400 2128.720 2663.000 2130.120 ;
        RECT 0.000 2113.800 2663.000 2128.720 ;
        RECT 0.000 2112.400 2662.600 2113.800 ;
        RECT 0.000 2104.280 2663.000 2112.400 ;
        RECT 0.000 2102.880 16.600 2104.280 ;
        RECT 21.400 2102.880 2663.000 2104.280 ;
        RECT 0.000 2087.960 2663.000 2102.880 ;
        RECT 0.000 2086.560 2662.600 2087.960 ;
        RECT 0.000 2079.800 2663.000 2086.560 ;
        RECT 0.000 2078.400 16.600 2079.800 ;
        RECT 21.400 2078.400 2663.000 2079.800 ;
        RECT 0.000 2063.480 2663.000 2078.400 ;
        RECT 0.000 2062.080 2662.600 2063.480 ;
        RECT 0.000 2055.320 2663.000 2062.080 ;
        RECT 0.000 2053.920 16.600 2055.320 ;
        RECT 21.400 2053.920 2663.000 2055.320 ;
        RECT 0.000 2039.000 2663.000 2053.920 ;
        RECT 0.000 2037.600 2662.600 2039.000 ;
        RECT 0.000 2030.840 2663.000 2037.600 ;
        RECT 0.000 2029.440 16.600 2030.840 ;
        RECT 21.400 2029.440 2663.000 2030.840 ;
        RECT 0.000 2014.520 2663.000 2029.440 ;
        RECT 0.000 2013.120 2662.600 2014.520 ;
        RECT 0.000 2005.000 2663.000 2013.120 ;
        RECT 0.000 2003.600 16.600 2005.000 ;
        RECT 21.400 2003.600 2663.000 2005.000 ;
        RECT 0.000 1990.040 2663.000 2003.600 ;
        RECT 0.000 1988.640 2662.600 1990.040 ;
        RECT 0.000 1980.520 2663.000 1988.640 ;
        RECT 0.000 1979.120 16.600 1980.520 ;
        RECT 21.400 1979.120 2663.000 1980.520 ;
        RECT 0.000 1964.200 2663.000 1979.120 ;
        RECT 0.000 1962.800 2662.600 1964.200 ;
        RECT 0.000 1956.040 2663.000 1962.800 ;
        RECT 0.000 1954.640 16.600 1956.040 ;
        RECT 21.400 1954.640 2663.000 1956.040 ;
        RECT 0.000 1939.720 2663.000 1954.640 ;
        RECT 0.000 1938.320 2662.600 1939.720 ;
        RECT 0.000 1931.560 2663.000 1938.320 ;
        RECT 0.000 1930.160 16.600 1931.560 ;
        RECT 21.400 1930.160 2663.000 1931.560 ;
        RECT 0.000 1915.240 2663.000 1930.160 ;
        RECT 0.000 1913.840 2662.600 1915.240 ;
        RECT 0.000 1905.720 2663.000 1913.840 ;
        RECT 0.000 1904.320 16.600 1905.720 ;
        RECT 21.400 1904.320 2663.000 1905.720 ;
        RECT 0.000 1890.760 2663.000 1904.320 ;
        RECT 0.000 1889.360 2662.600 1890.760 ;
        RECT 0.000 1881.240 2663.000 1889.360 ;
        RECT 0.000 1879.840 16.600 1881.240 ;
        RECT 21.400 1879.840 2663.000 1881.240 ;
        RECT 0.000 1864.920 2663.000 1879.840 ;
        RECT 0.000 1863.520 2662.600 1864.920 ;
        RECT 0.000 1856.760 2663.000 1863.520 ;
        RECT 0.000 1855.360 16.600 1856.760 ;
        RECT 21.400 1855.360 2663.000 1856.760 ;
        RECT 0.000 1840.440 2663.000 1855.360 ;
        RECT 0.000 1839.040 2662.600 1840.440 ;
        RECT 0.000 1832.280 2663.000 1839.040 ;
        RECT 0.000 1830.880 16.600 1832.280 ;
        RECT 21.400 1830.880 2663.000 1832.280 ;
        RECT 0.000 1815.960 2663.000 1830.880 ;
        RECT 0.000 1814.560 2662.600 1815.960 ;
        RECT 0.000 1807.800 2663.000 1814.560 ;
        RECT 0.000 1806.400 16.600 1807.800 ;
        RECT 21.400 1806.400 2663.000 1807.800 ;
        RECT 0.000 1791.480 2663.000 1806.400 ;
        RECT 0.000 1790.080 2662.600 1791.480 ;
        RECT 0.000 1781.960 2663.000 1790.080 ;
        RECT 0.000 1780.560 16.600 1781.960 ;
        RECT 21.400 1780.560 2663.000 1781.960 ;
        RECT 0.000 1765.640 2663.000 1780.560 ;
        RECT 0.000 1764.240 2662.600 1765.640 ;
        RECT 0.000 1757.480 2663.000 1764.240 ;
        RECT 0.000 1756.080 16.600 1757.480 ;
        RECT 21.400 1756.080 2663.000 1757.480 ;
        RECT 0.000 1741.160 2663.000 1756.080 ;
        RECT 0.000 1739.760 2662.600 1741.160 ;
        RECT 0.000 1733.000 2663.000 1739.760 ;
        RECT 0.000 1731.600 16.600 1733.000 ;
        RECT 21.400 1731.600 2663.000 1733.000 ;
        RECT 0.000 1716.680 2663.000 1731.600 ;
        RECT 0.000 1715.280 2662.600 1716.680 ;
        RECT 0.000 1708.520 2663.000 1715.280 ;
        RECT 0.000 1707.120 16.600 1708.520 ;
        RECT 21.400 1707.120 2663.000 1708.520 ;
        RECT 0.000 1692.200 2663.000 1707.120 ;
        RECT 0.000 1690.800 2662.600 1692.200 ;
        RECT 0.000 1682.680 2663.000 1690.800 ;
        RECT 0.000 1681.280 16.600 1682.680 ;
        RECT 21.400 1681.280 2663.000 1682.680 ;
        RECT 0.000 1666.360 2663.000 1681.280 ;
        RECT 0.000 1664.960 2662.600 1666.360 ;
        RECT 0.000 1658.200 2663.000 1664.960 ;
        RECT 0.000 1656.800 16.600 1658.200 ;
        RECT 21.400 1656.800 2663.000 1658.200 ;
        RECT 0.000 1641.880 2663.000 1656.800 ;
        RECT 0.000 1640.480 2662.600 1641.880 ;
        RECT 0.000 1633.720 2663.000 1640.480 ;
        RECT 0.000 1632.320 16.600 1633.720 ;
        RECT 21.400 1632.320 2663.000 1633.720 ;
        RECT 0.000 1617.400 2663.000 1632.320 ;
        RECT 0.000 1616.000 2662.600 1617.400 ;
        RECT 0.000 1609.240 2663.000 1616.000 ;
        RECT 0.000 1607.840 16.600 1609.240 ;
        RECT 21.400 1607.840 2663.000 1609.240 ;
        RECT 0.000 1592.920 2663.000 1607.840 ;
        RECT 0.000 1591.520 2662.600 1592.920 ;
        RECT 0.000 1583.400 2663.000 1591.520 ;
        RECT 0.000 1582.000 16.600 1583.400 ;
        RECT 21.400 1582.000 2663.000 1583.400 ;
        RECT 0.000 1568.440 2663.000 1582.000 ;
        RECT 0.000 1567.040 2662.600 1568.440 ;
        RECT 0.000 1558.920 2663.000 1567.040 ;
        RECT 0.000 1557.520 16.600 1558.920 ;
        RECT 21.400 1557.520 2663.000 1558.920 ;
        RECT 0.000 1542.600 2663.000 1557.520 ;
        RECT 0.000 1541.200 2662.600 1542.600 ;
        RECT 0.000 1534.440 2663.000 1541.200 ;
        RECT 0.000 1533.040 16.600 1534.440 ;
        RECT 21.400 1533.040 2663.000 1534.440 ;
        RECT 0.000 1518.120 2663.000 1533.040 ;
        RECT 0.000 1516.720 2662.600 1518.120 ;
        RECT 0.000 1509.960 2663.000 1516.720 ;
        RECT 0.000 1508.560 16.600 1509.960 ;
        RECT 21.400 1508.560 2663.000 1509.960 ;
        RECT 0.000 1493.640 2663.000 1508.560 ;
        RECT 0.000 1492.240 2662.600 1493.640 ;
        RECT 0.000 1484.120 2663.000 1492.240 ;
        RECT 0.000 1482.720 16.600 1484.120 ;
        RECT 21.400 1482.720 2663.000 1484.120 ;
        RECT 0.000 1469.160 2663.000 1482.720 ;
        RECT 0.000 1467.760 2662.600 1469.160 ;
        RECT 0.000 1459.640 2663.000 1467.760 ;
        RECT 0.000 1458.240 16.600 1459.640 ;
        RECT 21.400 1458.240 2663.000 1459.640 ;
        RECT 0.000 1443.320 2663.000 1458.240 ;
        RECT 0.000 1441.920 2662.600 1443.320 ;
        RECT 0.000 1435.160 2663.000 1441.920 ;
        RECT 0.000 1433.760 16.600 1435.160 ;
        RECT 21.400 1433.760 2663.000 1435.160 ;
        RECT 0.000 1418.840 2663.000 1433.760 ;
        RECT 0.000 1417.440 2662.600 1418.840 ;
        RECT 0.000 1410.680 2663.000 1417.440 ;
        RECT 0.000 1409.280 16.600 1410.680 ;
        RECT 21.400 1409.280 2663.000 1410.680 ;
        RECT 0.000 1394.360 2663.000 1409.280 ;
        RECT 0.000 1392.960 2662.600 1394.360 ;
        RECT 0.000 1386.200 2663.000 1392.960 ;
        RECT 0.000 1384.800 16.600 1386.200 ;
        RECT 21.400 1384.800 2663.000 1386.200 ;
        RECT 0.000 1369.880 2663.000 1384.800 ;
        RECT 0.000 1368.480 2662.600 1369.880 ;
        RECT 0.000 1360.360 2663.000 1368.480 ;
        RECT 0.000 1358.960 16.600 1360.360 ;
        RECT 21.400 1358.960 2663.000 1360.360 ;
        RECT 0.000 1344.040 2663.000 1358.960 ;
        RECT 0.000 1342.640 2662.600 1344.040 ;
        RECT 0.000 1335.880 2663.000 1342.640 ;
        RECT 0.000 1334.480 16.600 1335.880 ;
        RECT 21.400 1334.480 2663.000 1335.880 ;
        RECT 0.000 1319.560 2663.000 1334.480 ;
        RECT 0.000 1318.160 2662.600 1319.560 ;
        RECT 0.000 1311.400 2663.000 1318.160 ;
        RECT 0.000 1310.000 16.600 1311.400 ;
        RECT 21.400 1310.000 2663.000 1311.400 ;
        RECT 0.000 1295.080 2663.000 1310.000 ;
        RECT 0.000 1293.680 2662.600 1295.080 ;
        RECT 0.000 1286.920 2663.000 1293.680 ;
        RECT 0.000 1285.520 16.600 1286.920 ;
        RECT 21.400 1285.520 2663.000 1286.920 ;
        RECT 0.000 1270.600 2663.000 1285.520 ;
        RECT 0.000 1269.200 2662.600 1270.600 ;
        RECT 0.000 1261.080 2663.000 1269.200 ;
        RECT 0.000 1259.680 16.600 1261.080 ;
        RECT 21.400 1259.680 2663.000 1261.080 ;
        RECT 0.000 1244.760 2663.000 1259.680 ;
        RECT 0.000 1243.360 2662.600 1244.760 ;
        RECT 0.000 1236.600 2663.000 1243.360 ;
        RECT 0.000 1235.200 16.600 1236.600 ;
        RECT 21.400 1235.200 2663.000 1236.600 ;
        RECT 0.000 1220.280 2663.000 1235.200 ;
        RECT 0.000 1218.880 2662.600 1220.280 ;
        RECT 0.000 1212.120 2663.000 1218.880 ;
        RECT 0.000 1210.720 16.600 1212.120 ;
        RECT 21.400 1210.720 2663.000 1212.120 ;
        RECT 0.000 1195.800 2663.000 1210.720 ;
        RECT 0.000 1194.400 2662.600 1195.800 ;
        RECT 0.000 1187.640 2663.000 1194.400 ;
        RECT 0.000 1186.240 16.600 1187.640 ;
        RECT 21.400 1186.240 2663.000 1187.640 ;
        RECT 0.000 1171.320 2663.000 1186.240 ;
        RECT 0.000 1169.920 2662.600 1171.320 ;
        RECT 0.000 1161.800 2663.000 1169.920 ;
        RECT 0.000 1160.400 16.600 1161.800 ;
        RECT 21.400 1160.400 2663.000 1161.800 ;
        RECT 0.000 1146.840 2663.000 1160.400 ;
        RECT 0.000 1145.440 2662.600 1146.840 ;
        RECT 0.000 1137.320 2663.000 1145.440 ;
        RECT 0.000 1135.920 16.600 1137.320 ;
        RECT 21.400 1135.920 2663.000 1137.320 ;
        RECT 0.000 1121.000 2663.000 1135.920 ;
        RECT 0.000 1119.600 2662.600 1121.000 ;
        RECT 0.000 1112.840 2663.000 1119.600 ;
        RECT 0.000 1111.440 16.600 1112.840 ;
        RECT 21.400 1111.440 2663.000 1112.840 ;
        RECT 0.000 1096.520 2663.000 1111.440 ;
        RECT 0.000 1095.120 2662.600 1096.520 ;
        RECT 0.000 1088.360 2663.000 1095.120 ;
        RECT 0.000 1086.960 16.600 1088.360 ;
        RECT 21.400 1086.960 2663.000 1088.360 ;
        RECT 0.000 1072.040 2663.000 1086.960 ;
        RECT 0.000 1070.640 2662.600 1072.040 ;
        RECT 0.000 1062.520 2663.000 1070.640 ;
        RECT 0.000 1061.120 16.600 1062.520 ;
        RECT 21.400 1061.120 2663.000 1062.520 ;
        RECT 0.000 1047.560 2663.000 1061.120 ;
        RECT 0.000 1046.160 2662.600 1047.560 ;
        RECT 0.000 1038.040 2663.000 1046.160 ;
        RECT 0.000 1036.640 16.600 1038.040 ;
        RECT 21.400 1036.640 2663.000 1038.040 ;
        RECT 0.000 1021.720 2663.000 1036.640 ;
        RECT 0.000 1020.320 2662.600 1021.720 ;
        RECT 0.000 1013.560 2663.000 1020.320 ;
        RECT 0.000 1012.160 16.600 1013.560 ;
        RECT 21.400 1012.160 2663.000 1013.560 ;
        RECT 0.000 997.240 2663.000 1012.160 ;
        RECT 0.000 995.840 2662.600 997.240 ;
        RECT 0.000 989.080 2663.000 995.840 ;
        RECT 0.000 987.680 16.600 989.080 ;
        RECT 21.400 987.680 2663.000 989.080 ;
        RECT 0.000 972.760 2663.000 987.680 ;
        RECT 0.000 971.360 2662.600 972.760 ;
        RECT 0.000 963.240 2663.000 971.360 ;
        RECT 0.000 961.840 16.600 963.240 ;
        RECT 21.400 961.840 2663.000 963.240 ;
        RECT 0.000 948.280 2663.000 961.840 ;
        RECT 0.000 946.880 2662.600 948.280 ;
        RECT 0.000 938.760 2663.000 946.880 ;
        RECT 0.000 937.360 16.600 938.760 ;
        RECT 21.400 937.360 2663.000 938.760 ;
        RECT 0.000 922.440 2663.000 937.360 ;
        RECT 0.000 921.040 2662.600 922.440 ;
        RECT 0.000 914.280 2663.000 921.040 ;
        RECT 0.000 912.880 16.600 914.280 ;
        RECT 21.400 912.880 2663.000 914.280 ;
        RECT 0.000 897.960 2663.000 912.880 ;
        RECT 0.000 896.560 2662.600 897.960 ;
        RECT 0.000 889.800 2663.000 896.560 ;
        RECT 0.000 888.400 16.600 889.800 ;
        RECT 21.400 888.400 2663.000 889.800 ;
        RECT 0.000 873.480 2663.000 888.400 ;
        RECT 0.000 872.080 2662.600 873.480 ;
        RECT 0.000 865.320 2663.000 872.080 ;
        RECT 0.000 863.920 16.600 865.320 ;
        RECT 21.400 863.920 2663.000 865.320 ;
        RECT 0.000 849.000 2663.000 863.920 ;
        RECT 0.000 847.600 2662.600 849.000 ;
        RECT 0.000 839.480 2663.000 847.600 ;
        RECT 0.000 838.080 16.600 839.480 ;
        RECT 21.400 838.080 2663.000 839.480 ;
        RECT 0.000 823.160 2663.000 838.080 ;
        RECT 0.000 821.760 2662.600 823.160 ;
        RECT 0.000 815.000 2663.000 821.760 ;
        RECT 0.000 813.600 16.600 815.000 ;
        RECT 21.400 813.600 2663.000 815.000 ;
        RECT 0.000 798.680 2663.000 813.600 ;
        RECT 0.000 797.280 2662.600 798.680 ;
        RECT 0.000 790.520 2663.000 797.280 ;
        RECT 0.000 789.120 16.600 790.520 ;
        RECT 21.400 789.120 2663.000 790.520 ;
        RECT 0.000 774.200 2663.000 789.120 ;
        RECT 0.000 772.800 2662.600 774.200 ;
        RECT 0.000 766.040 2663.000 772.800 ;
        RECT 0.000 764.640 16.600 766.040 ;
        RECT 21.400 764.640 2663.000 766.040 ;
        RECT 0.000 749.720 2663.000 764.640 ;
        RECT 0.000 748.320 2662.600 749.720 ;
        RECT 0.000 740.200 2663.000 748.320 ;
        RECT 0.000 738.800 16.600 740.200 ;
        RECT 21.400 738.800 2663.000 740.200 ;
        RECT 0.000 723.880 2663.000 738.800 ;
        RECT 0.000 722.480 2662.600 723.880 ;
        RECT 0.000 715.720 2663.000 722.480 ;
        RECT 0.000 714.320 16.600 715.720 ;
        RECT 21.400 714.320 2663.000 715.720 ;
        RECT 0.000 699.400 2663.000 714.320 ;
        RECT 0.000 698.000 2662.600 699.400 ;
        RECT 0.000 691.240 2663.000 698.000 ;
        RECT 0.000 689.840 16.600 691.240 ;
        RECT 21.400 689.840 2663.000 691.240 ;
        RECT 0.000 674.920 2663.000 689.840 ;
        RECT 0.000 673.520 2662.600 674.920 ;
        RECT 0.000 666.760 2663.000 673.520 ;
        RECT 0.000 665.360 16.600 666.760 ;
        RECT 21.400 665.360 2663.000 666.760 ;
        RECT 0.000 650.440 2663.000 665.360 ;
        RECT 0.000 649.040 2662.600 650.440 ;
        RECT 0.000 640.920 2663.000 649.040 ;
        RECT 0.000 639.520 16.600 640.920 ;
        RECT 21.400 639.520 2663.000 640.920 ;
        RECT 0.000 625.960 2663.000 639.520 ;
        RECT 0.000 624.560 2662.600 625.960 ;
        RECT 0.000 616.440 2663.000 624.560 ;
        RECT 0.000 615.040 16.600 616.440 ;
        RECT 21.400 615.040 2663.000 616.440 ;
        RECT 0.000 600.120 2663.000 615.040 ;
        RECT 0.000 598.720 2662.600 600.120 ;
        RECT 0.000 591.960 2663.000 598.720 ;
        RECT 0.000 590.560 16.600 591.960 ;
        RECT 21.400 590.560 2663.000 591.960 ;
        RECT 0.000 575.640 2663.000 590.560 ;
        RECT 0.000 574.240 2662.600 575.640 ;
        RECT 0.000 567.480 2663.000 574.240 ;
        RECT 0.000 566.080 16.600 567.480 ;
        RECT 21.400 566.080 2663.000 567.480 ;
        RECT 0.000 551.160 2663.000 566.080 ;
        RECT 0.000 549.760 2662.600 551.160 ;
        RECT 0.000 541.640 2663.000 549.760 ;
        RECT 0.000 540.240 16.600 541.640 ;
        RECT 21.400 540.240 2663.000 541.640 ;
        RECT 0.000 526.680 2663.000 540.240 ;
        RECT 0.000 525.280 2662.600 526.680 ;
        RECT 0.000 517.160 2663.000 525.280 ;
        RECT 0.000 515.760 16.600 517.160 ;
        RECT 21.400 515.760 2663.000 517.160 ;
        RECT 0.000 500.840 2663.000 515.760 ;
        RECT 0.000 499.440 2662.600 500.840 ;
        RECT 0.000 492.680 2663.000 499.440 ;
        RECT 0.000 491.280 16.600 492.680 ;
        RECT 21.400 491.280 2663.000 492.680 ;
        RECT 0.000 476.360 2663.000 491.280 ;
        RECT 0.000 474.960 2662.600 476.360 ;
        RECT 0.000 468.200 2663.000 474.960 ;
        RECT 0.000 466.800 16.600 468.200 ;
        RECT 21.400 466.800 2663.000 468.200 ;
        RECT 0.000 451.880 2663.000 466.800 ;
        RECT 0.000 450.480 2662.600 451.880 ;
        RECT 0.000 443.720 2663.000 450.480 ;
        RECT 0.000 442.320 16.600 443.720 ;
        RECT 21.400 442.320 2663.000 443.720 ;
        RECT 0.000 427.400 2663.000 442.320 ;
        RECT 0.000 426.000 2662.600 427.400 ;
        RECT 0.000 417.880 2663.000 426.000 ;
        RECT 0.000 416.480 16.600 417.880 ;
        RECT 21.400 416.480 2663.000 417.880 ;
        RECT 0.000 401.560 2663.000 416.480 ;
        RECT 0.000 400.160 2662.600 401.560 ;
        RECT 0.000 393.400 2663.000 400.160 ;
        RECT 0.000 392.000 16.600 393.400 ;
        RECT 21.400 392.000 2663.000 393.400 ;
        RECT 0.000 377.080 2663.000 392.000 ;
        RECT 0.000 375.680 2662.600 377.080 ;
        RECT 0.000 368.920 2663.000 375.680 ;
        RECT 0.000 367.520 16.600 368.920 ;
        RECT 21.400 367.520 2663.000 368.920 ;
        RECT 0.000 352.600 2663.000 367.520 ;
        RECT 0.000 351.200 2662.600 352.600 ;
        RECT 0.000 344.440 2663.000 351.200 ;
        RECT 0.000 343.040 16.600 344.440 ;
        RECT 21.400 343.040 2663.000 344.440 ;
        RECT 0.000 328.120 2663.000 343.040 ;
        RECT 0.000 326.720 2662.600 328.120 ;
        RECT 0.000 318.600 2663.000 326.720 ;
        RECT 0.000 317.200 16.600 318.600 ;
        RECT 21.400 317.200 2663.000 318.600 ;
        RECT 0.000 302.280 2663.000 317.200 ;
        RECT 0.000 300.880 2662.600 302.280 ;
        RECT 0.000 294.120 2663.000 300.880 ;
        RECT 0.000 292.720 16.600 294.120 ;
        RECT 21.400 292.720 2663.000 294.120 ;
        RECT 0.000 277.800 2663.000 292.720 ;
        RECT 0.000 276.400 2662.600 277.800 ;
        RECT 0.000 269.640 2663.000 276.400 ;
        RECT 0.000 268.240 16.600 269.640 ;
        RECT 21.400 268.240 2663.000 269.640 ;
        RECT 0.000 253.320 2663.000 268.240 ;
        RECT 0.000 251.920 2662.600 253.320 ;
        RECT 0.000 245.160 2663.000 251.920 ;
        RECT 0.000 243.760 16.600 245.160 ;
        RECT 21.400 243.760 2663.000 245.160 ;
        RECT 0.000 228.840 2663.000 243.760 ;
        RECT 0.000 227.440 2662.600 228.840 ;
        RECT 0.000 219.320 2663.000 227.440 ;
        RECT 0.000 217.920 16.600 219.320 ;
        RECT 21.400 217.920 2663.000 219.320 ;
        RECT 0.000 204.360 2663.000 217.920 ;
        RECT 0.000 202.960 2662.600 204.360 ;
        RECT 0.000 194.840 2663.000 202.960 ;
        RECT 0.000 193.440 16.600 194.840 ;
        RECT 21.400 193.440 2663.000 194.840 ;
        RECT 0.000 178.520 2663.000 193.440 ;
        RECT 0.000 177.120 2662.600 178.520 ;
        RECT 0.000 170.360 2663.000 177.120 ;
        RECT 0.000 168.960 16.600 170.360 ;
        RECT 21.400 168.960 2663.000 170.360 ;
        RECT 0.000 154.040 2663.000 168.960 ;
        RECT 0.000 152.640 2662.600 154.040 ;
        RECT 0.000 145.880 2663.000 152.640 ;
        RECT 0.000 144.480 16.600 145.880 ;
        RECT 21.400 144.480 2663.000 145.880 ;
        RECT 0.000 129.560 2663.000 144.480 ;
        RECT 0.000 128.160 2662.600 129.560 ;
        RECT 0.000 120.040 2663.000 128.160 ;
        RECT 0.000 118.640 16.600 120.040 ;
        RECT 21.400 118.640 2663.000 120.040 ;
        RECT 0.000 105.080 2663.000 118.640 ;
        RECT 0.000 103.680 2662.600 105.080 ;
        RECT 0.000 95.560 2663.000 103.680 ;
        RECT 0.000 94.160 16.600 95.560 ;
        RECT 21.400 94.160 2663.000 95.560 ;
        RECT 0.000 79.240 2663.000 94.160 ;
        RECT 0.000 77.840 2662.600 79.240 ;
        RECT 0.000 71.080 2663.000 77.840 ;
        RECT 0.000 69.680 16.600 71.080 ;
        RECT 21.400 69.680 2663.000 71.080 ;
        RECT 0.000 54.760 2663.000 69.680 ;
        RECT 0.000 53.360 2662.600 54.760 ;
        RECT 0.000 46.600 2663.000 53.360 ;
        RECT 0.000 45.200 16.600 46.600 ;
        RECT 21.400 45.200 2663.000 46.600 ;
        RECT 0.000 30.280 2663.000 45.200 ;
        RECT 0.000 28.880 2662.600 30.280 ;
        RECT 0.000 0.000 2663.000 28.880 ;
      LAYER met4 ;
        RECT 22.815 16.760 2653.425 3645.985 ;
      LAYER met5 ;
        RECT 17.000 185.790 2623.480 3643.900 ;
  END
END ghazi_top_dffram_csv
END LIBRARY

