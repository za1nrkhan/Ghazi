VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ghazi_top_dffram_csv
  CLASS BLOCK ;
  FOREIGN ghazi_top_dffram_csv ;
  ORIGIN 0.000 0.000 ;
  SIZE 2700.000 BY 3470.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.290 3466.000 9.570 3470.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1521.880 2700.000 1522.480 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2043.410 3466.000 2043.690 3470.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.570 0.000 2202.850 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1788.440 4.000 1789.040 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.890 3466.000 175.170 3470.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1514.410 3466.000 1514.690 3470.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2632.210 0.000 2632.490 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1050.730 3466.000 1051.010 3470.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1032.280 2700.000 1032.880 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1347.800 4.000 1348.400 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1993.730 3466.000 1994.010 3470.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 250.280 2700.000 250.880 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1006.440 4.000 1007.040 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1396.760 4.000 1397.360 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2769.000 2700.000 2769.600 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 647.770 0.000 648.050 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3084.520 4.000 3085.120 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2582.530 0.000 2582.810 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1034.170 3466.000 1034.450 3470.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1166.650 3466.000 1166.930 3470.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 968.850 3466.000 969.130 3470.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.930 0.000 1359.210 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2842.440 2700.000 2843.040 ;
    END
  END io_in[36]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.890 3466.000 2590.170 3470.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2084.920 2700.000 2085.520 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1093.970 0.000 1094.250 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3405.480 2700.000 3406.080 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1464.730 3466.000 1465.010 3470.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.650 3466.000 108.930 3470.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 472.050 3466.000 472.330 3470.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2060.440 2700.000 2061.040 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3111.720 2700.000 3112.320 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1717.720 2700.000 1718.320 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 908.520 4.000 909.120 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 505.170 3466.000 505.450 3470.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 617.480 2700.000 618.080 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 4.000 737.760 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1668.760 2700.000 1669.360 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2136.330 0.000 2136.610 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 621.090 3466.000 621.370 3470.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3062.760 2700.000 3063.360 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1877.810 3466.000 1878.090 3470.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1644.280 2700.000 1644.880 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.720 4.000 1446.320 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2219.130 0.000 2219.410 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1772.010 0.000 1772.290 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3454.440 2700.000 3455.040 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2407.730 3466.000 2408.010 3470.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2665.330 0.000 2665.610 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1398.490 3466.000 1398.770 3470.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1372.280 4.000 1372.880 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1607.330 0.000 1607.610 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 3466.000 92.370 3470.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3231.400 4.000 3232.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1568.120 4.000 1568.720 ;
    END
  END io_oeb[36]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3402.760 4.000 3403.360 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2182.840 2700.000 2183.440 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2540.210 3466.000 2540.490 3470.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 720.450 3466.000 720.730 3470.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.690 3466.000 2672.970 3470.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1408.610 0.000 1408.890 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2142.770 3466.000 2143.050 3470.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 554.850 3466.000 555.130 3470.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 422.370 3466.000 422.650 3470.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 730.570 0.000 730.850 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2053.530 0.000 2053.810 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2152.890 0.000 2153.170 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1987.000 2700.000 1987.600 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3185.160 2700.000 3185.760 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2790.760 4.000 2791.360 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1580.650 3466.000 1580.930 3470.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.720 4.000 664.320 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1657.010 0.000 1657.290 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2401.290 0.000 2401.570 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2254.920 2700.000 2255.520 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2400.440 4.000 2401.040 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 571.410 3466.000 571.690 3470.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1592.600 4.000 1593.200 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3307.560 2700.000 3308.160 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1133.530 3466.000 1133.810 3470.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 862.280 2700.000 862.880 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1646.890 3466.000 1647.170 3470.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1017.610 3466.000 1017.890 3470.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 339.570 3466.000 339.850 3470.000 ;
    END
  END io_out[36]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1007.800 2700.000 1008.400 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1910.840 4.000 1911.440 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3258.600 2700.000 3259.200 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1696.570 3466.000 1696.850 3470.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1399.480 2700.000 1400.080 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1763.960 4.000 1764.560 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2209.010 3466.000 2209.290 3470.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1640.450 0.000 1640.730 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.530 3466.000 190.810 3470.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1425.170 0.000 1425.450 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 788.840 2700.000 789.440 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 323.720 2700.000 324.320 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 737.010 3466.000 737.290 3470.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2358.050 3466.000 2358.330 3470.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1746.250 3466.000 1746.530 3470.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2301.930 0.000 2302.210 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1323.320 4.000 1323.920 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1203.640 2700.000 1204.240 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.650 3466.000 2523.930 3470.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2327.000 4.000 2327.600 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1104.360 4.000 1104.960 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2450.970 0.000 2451.250 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2615.650 0.000 2615.930 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 770.130 3466.000 770.410 3470.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1177.800 4.000 1178.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1960.610 3466.000 1960.890 3470.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1887.930 0.000 1888.210 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3255.880 4.000 3256.480 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 859.560 4.000 860.160 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2619.400 4.000 2620.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2497.000 4.000 2497.600 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1595.320 2700.000 1595.920 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.000 4.000 933.600 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 201.320 2700.000 201.920 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2744.520 2700.000 2745.120 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3378.280 4.000 3378.880 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2689.250 3466.000 2689.530 3470.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 952.290 3466.000 952.570 3470.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 521.730 3466.000 522.010 3470.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2681.890 0.000 2682.170 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2192.450 3466.000 2192.730 3470.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 984.680 2700.000 985.280 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1921.050 0.000 1921.330 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3209.640 2700.000 3210.240 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1913.560 2700.000 1914.160 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2401.800 2700.000 2402.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 803.250 3466.000 803.530 3470.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1959.800 4.000 1960.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 960.200 2700.000 960.800 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 687.330 3466.000 687.610 3470.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2204.600 4.000 2205.200 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3283.080 2700.000 3283.680 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1619.800 2700.000 1620.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2695.560 2700.000 2696.160 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1829.050 3466.000 1829.330 3470.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2594.920 4.000 2595.520 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3011.080 4.000 3011.680 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2915.880 2700.000 2916.480 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2548.680 2700.000 2549.280 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2668.360 4.000 2668.960 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1597.210 3466.000 1597.490 3470.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2962.120 4.000 2962.720 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 886.760 2700.000 887.360 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1630.330 3466.000 1630.610 3470.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3206.920 4.000 3207.520 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 911.810 0.000 912.090 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2335.050 0.000 2335.330 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1861.250 3466.000 1861.530 3470.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2622.120 2700.000 2622.720 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1202.280 4.000 1202.880 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1864.600 2700.000 1865.200 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1944.050 3466.000 1944.330 3470.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2556.770 3466.000 2557.050 3470.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3136.200 2700.000 3136.800 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3234.120 2700.000 3234.720 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.210 0.000 2517.490 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 127.880 2700.000 128.480 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2103.210 0.000 2103.490 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1079.880 4.000 1080.480 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2010.290 3466.000 2010.570 3470.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 421.640 2700.000 422.240 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1984.280 4.000 1984.880 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1927.490 3466.000 1927.770 3470.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1871.370 0.000 1871.650 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1546.360 2700.000 1546.960 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3035.560 4.000 3036.160 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2449.400 4.000 2450.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3356.520 2700.000 3357.120 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1613.770 3466.000 1614.050 3470.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2351.610 0.000 2351.890 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1519.160 4.000 1519.760 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.410 3466.000 42.690 3470.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.250 3466.000 389.530 3470.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1350.520 2700.000 1351.120 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 593.000 2700.000 593.600 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1055.400 4.000 1056.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2599.090 0.000 2599.370 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2158.360 2700.000 2158.960 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2318.490 0.000 2318.770 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 225.800 2700.000 226.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3160.680 2700.000 3161.280 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.090 3466.000 1150.370 3470.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1689.210 0.000 1689.490 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2815.240 4.000 2815.840 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 981.960 4.000 982.560 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2285.370 0.000 2285.650 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 538.290 3466.000 538.570 3470.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 78.920 2700.000 79.520 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 902.610 3466.000 902.890 3470.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2275.250 3466.000 2275.530 3470.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1739.480 4.000 1740.080 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1160.210 0.000 1160.490 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.690 3466.000 372.970 3470.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 935.720 2700.000 936.320 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2570.440 4.000 2571.040 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2020.410 0.000 2020.690 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2230.440 2700.000 2231.040 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1861.880 4.000 1862.480 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1392.050 0.000 1392.330 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2648.770 0.000 2649.050 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 372.680 2700.000 373.280 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1791.160 2700.000 1791.760 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 928.370 0.000 928.650 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2839.720 4.000 2840.320 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2741.800 4.000 2742.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2643.880 4.000 2644.480 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2473.970 3466.000 2474.250 3470.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1507.970 0.000 1508.250 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3304.840 4.000 3305.440 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1755.450 0.000 1755.730 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2008.760 4.000 2009.360 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2341.490 3466.000 2341.770 3470.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3332.040 2700.000 3332.640 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2003.850 0.000 2004.130 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1375.000 2700.000 1375.600 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1766.680 2700.000 1767.280 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2229.080 4.000 2229.680 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 935.730 3466.000 936.010 3470.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 240.210 3466.000 240.490 3470.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 957.480 4.000 958.080 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 944.930 0.000 945.210 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1795.930 3466.000 1796.210 3470.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 911.240 2700.000 911.840 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.730 0.000 1442.010 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2467.530 0.000 2467.810 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1481.290 3466.000 1481.570 3470.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1729.690 3466.000 1729.970 3470.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1143.650 0.000 1143.930 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 5.480 2700.000 6.080 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 604.530 3466.000 604.810 3470.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.770 0.000 2120.050 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2671.080 2700.000 2671.680 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1266.010 3466.000 1266.290 3470.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2964.840 2700.000 2965.440 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 637.650 3466.000 637.930 3470.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2131.160 4.000 2131.760 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1252.600 2700.000 1253.200 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1543.640 4.000 1544.240 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3087.240 2700.000 3087.840 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2109.400 2700.000 2110.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2155.640 4.000 2156.240 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1497.400 2700.000 1498.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 498.730 0.000 499.010 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1472.920 2700.000 1473.520 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2180.120 4.000 2180.720 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.170 3466.000 1977.450 3470.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 299.240 2700.000 299.840 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1056.760 2700.000 1057.360 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 715.400 2700.000 716.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1491.410 0.000 1491.690 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2499.720 2700.000 2500.320 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 158.330 3466.000 158.610 3470.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3182.440 4.000 3183.040 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1176.770 0.000 1177.050 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2076.530 3466.000 2076.810 3470.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1894.370 3466.000 1894.650 3470.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2133.880 2700.000 2134.480 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 836.370 3466.000 836.650 3470.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 961.490 0.000 961.770 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1298.840 4.000 1299.440 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1282.570 3466.000 1282.850 3470.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2639.570 3466.000 2639.850 3470.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 273.330 3466.000 273.610 3470.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1474.850 0.000 1475.130 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1274.360 4.000 1274.960 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2913.160 4.000 2913.760 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.890 0.000 1210.170 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2891.400 2700.000 2892.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2225.570 3466.000 2225.850 3470.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1680.010 3466.000 1680.290 3470.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1301.560 2700.000 1302.160 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1325.810 0.000 1326.090 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 4.000 713.280 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2720.040 2700.000 2720.640 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 54.440 2700.000 55.040 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1547.530 3466.000 1547.810 3470.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1840.120 2700.000 1840.720 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 813.370 0.000 813.650 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2026.850 3466.000 2027.130 3470.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1937.610 0.000 1937.890 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 994.610 0.000 994.890 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.290 0.000 1987.570 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2252.250 0.000 2252.530 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1216.330 3466.000 1216.610 3470.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1889.080 2700.000 1889.680 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2532.850 0.000 2533.130 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 446.120 2700.000 446.720 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 29.960 2700.000 30.560 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.690 3466.000 786.970 3470.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2573.330 3466.000 2573.610 3470.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1226.450 0.000 1226.730 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2368.170 0.000 2368.450 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1105.720 2700.000 1106.320 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 978.050 0.000 978.330 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1821.690 0.000 1821.970 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2126.210 3466.000 2126.490 3470.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1690.520 4.000 1691.120 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1962.520 2700.000 1963.120 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1854.810 0.000 1855.090 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2521.480 4.000 2522.080 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2070.090 0.000 2070.370 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2986.600 4.000 2987.200 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3133.480 4.000 3134.080 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1742.200 2700.000 1742.800 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.930 3466.000 853.210 3470.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1693.240 2700.000 1693.840 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 103.400 2700.000 104.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 256.770 3466.000 257.050 3470.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2490.530 3466.000 2490.810 3470.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2391.170 3466.000 2391.450 3470.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3329.320 4.000 3329.920 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2473.880 4.000 2474.480 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2646.600 2700.000 2647.200 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1249.450 3466.000 1249.730 3470.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1027.730 0.000 1028.010 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.530 0.000 1110.810 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2035.960 2700.000 2036.560 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1570.840 2700.000 1571.440 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1276.130 0.000 1276.410 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2793.480 2700.000 2794.080 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1100.410 3466.000 1100.690 3470.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2303.880 2700.000 2304.480 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1116.970 3466.000 1117.250 3470.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.610 3466.000 1845.890 3470.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1954.170 0.000 1954.450 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1342.370 0.000 1342.650 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2937.640 4.000 2938.240 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 753.570 3466.000 753.850 3470.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1381.930 3466.000 1382.210 3470.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1130.200 2700.000 1130.800 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1153.320 4.000 1153.920 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.970 3466.000 588.250 3470.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1762.810 3466.000 1763.090 3470.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 495.080 2700.000 495.680 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1348.810 3466.000 1349.090 3470.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 176.840 2700.000 177.440 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3381.000 2700.000 3381.600 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 739.880 2700.000 740.480 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1249.880 4.000 1250.480 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2159.330 3466.000 2159.610 3470.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.850 0.000 2418.130 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1154.680 2700.000 1155.280 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1277.080 2700.000 1277.680 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2597.640 2700.000 2598.240 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1497.850 3466.000 1498.130 3470.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1886.360 4.000 1886.960 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1292.690 0.000 1292.970 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1938.040 2700.000 1938.640 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1448.170 3466.000 1448.450 3470.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 837.800 2700.000 838.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2424.920 4.000 2425.520 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2475.240 2700.000 2475.840 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1259.570 0.000 1259.850 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.930 0.000 830.210 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 397.160 2700.000 397.760 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.530 0.000 1524.810 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 666.440 2700.000 667.040 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1541.090 0.000 1541.370 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.970 0.000 2037.250 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2549.410 0.000 2549.690 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 274.760 2700.000 275.360 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.490 3466.000 455.770 3470.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 223.650 3466.000 223.930 3470.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3353.800 4.000 3354.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2302.520 4.000 2303.120 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1641.560 4.000 1642.160 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2524.200 2700.000 2524.800 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2989.320 2700.000 2989.920 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2324.930 3466.000 2325.210 3470.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2573.160 2700.000 2573.760 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3109.000 4.000 3109.600 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 544.040 2700.000 544.640 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2242.130 3466.000 2242.410 3470.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2377.320 2700.000 2377.920 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1326.040 2700.000 1326.640 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1332.250 3466.000 1332.530 3470.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1530.970 3466.000 1531.250 3470.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 869.490 3466.000 869.770 3470.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2175.890 3466.000 2176.170 3470.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1375.490 0.000 1375.770 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2207.320 2700.000 2207.920 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 356.130 3466.000 356.410 3470.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2606.450 3466.000 2606.730 3470.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 306.450 3466.000 306.730 3470.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1910.930 3466.000 1911.210 3470.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2692.840 4.000 2693.440 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1421.240 4.000 1421.840 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2866.920 2700.000 2867.520 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 405.810 3466.000 406.090 3470.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2717.320 4.000 2717.920 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1199.770 3466.000 1200.050 3470.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.770 0.000 1591.050 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1448.440 2700.000 1449.040 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2235.690 0.000 2235.970 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.890 0.000 681.170 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2374.610 3466.000 2374.890 3470.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2033.240 4.000 2033.840 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1837.400 4.000 1838.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3038.280 2700.000 3038.880 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.080 4.000 835.680 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2766.280 4.000 2766.880 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1812.490 3466.000 1812.770 3470.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2291.810 3466.000 2292.090 3470.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2888.680 4.000 2889.280 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1179.160 2700.000 1179.760 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 862.130 0.000 862.410 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1243.010 0.000 1243.290 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 488.610 3466.000 488.890 3470.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1315.690 3466.000 1315.970 3470.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2352.840 2700.000 2353.440 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 289.890 3466.000 290.170 3470.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2864.200 4.000 2864.800 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3427.240 4.000 3427.840 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 813.320 2700.000 813.920 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1564.090 3466.000 1564.370 3470.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1228.120 2700.000 1228.720 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2817.960 2700.000 2818.560 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2623.010 3466.000 2623.290 3470.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 568.520 2700.000 569.120 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2253.560 4.000 2254.160 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 470.600 2700.000 471.200 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 985.410 3466.000 985.690 3470.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 690.920 2700.000 691.520 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1494.680 4.000 1495.280 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2093.090 3466.000 2093.370 3470.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.650 0.000 2500.930 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1713.130 3466.000 1713.410 3470.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.410 0.000 2434.690 4.000 ;
    END
  END la_oen[9]
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 348.200 2700.000 348.800 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2082.200 4.000 2082.800 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1970.730 0.000 1971.010 4.000 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1077.410 0.000 1077.690 4.000 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3157.960 4.000 3158.560 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1001.970 3466.000 1002.250 3470.000 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1617.080 4.000 1617.680 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3013.800 2700.000 3014.400 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1673.570 0.000 1673.850 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 664.330 0.000 664.610 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1788.570 0.000 1788.850 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 125.210 3466.000 125.490 3470.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3280.360 4.000 3280.960 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1365.370 3466.000 1365.650 3470.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 3466.000 26.130 3470.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2424.290 3466.000 2424.570 3470.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1779.370 3466.000 1779.650 3470.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1081.240 2700.000 1081.840 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1011.170 0.000 1011.450 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1470.200 4.000 1470.800 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1812.920 4.000 1813.520 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1226.760 4.000 1227.360 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1232.890 3466.000 1233.170 3470.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2507.090 3466.000 2507.370 3470.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1935.320 4.000 1935.920 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 519.560 2700.000 520.160 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2450.760 2700.000 2451.360 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1183.210 3466.000 1183.490 3470.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 670.770 3466.000 671.050 3470.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2426.280 2700.000 2426.880 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2086.650 0.000 2086.930 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 845.570 0.000 845.850 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1044.290 0.000 1044.570 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1299.130 3466.000 1299.410 3470.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2384.730 0.000 2385.010 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1423.960 2700.000 1424.560 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1838.250 0.000 1838.530 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.850 3466.000 1084.130 3470.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1557.650 0.000 1557.930 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1805.130 0.000 1805.410 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 810.600 4.000 811.200 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2186.010 0.000 2186.290 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 207.090 3466.000 207.370 3470.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1309.250 0.000 1309.530 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1715.000 4.000 1715.600 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2457.410 3466.000 2457.690 3470.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2440.850 3466.000 2441.130 3470.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3429.960 2700.000 3430.560 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2109.650 3466.000 2109.930 3470.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1060.850 0.000 1061.130 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.770 3466.000 142.050 3470.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2545.960 4.000 2546.560 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1415.050 3466.000 1415.330 3470.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2279.400 2700.000 2280.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2328.360 2700.000 2328.960 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 3466.000 59.250 3470.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 878.690 0.000 878.970 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 641.960 2700.000 642.560 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 764.360 2700.000 764.960 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.810 0.000 2269.090 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2011.480 2700.000 2012.080 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1705.770 0.000 1706.050 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1193.330 0.000 1193.610 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1722.330 0.000 1722.610 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2375.960 4.000 2376.560 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2484.090 0.000 2484.370 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1431.610 3466.000 1431.890 3470.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 919.170 3466.000 919.450 3470.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2258.690 3466.000 2258.970 3470.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2057.720 4.000 2058.320 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.290 3466.000 1067.570 3470.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.970 0.000 2566.250 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1666.040 4.000 1666.640 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 152.360 2700.000 152.960 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1458.290 0.000 1458.570 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.920 4.000 1031.520 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.530 3466.000 75.810 3470.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2656.130 3466.000 2656.410 3470.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1623.890 0.000 1624.170 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2308.370 3466.000 2308.650 3470.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.930 3466.000 439.210 3470.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 819.810 3466.000 820.090 3470.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1904.490 0.000 1904.770 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2169.450 0.000 2169.730 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2278.040 4.000 2278.640 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 654.210 3466.000 654.490 3470.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2351.480 4.000 2352.080 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2940.360 2700.000 2940.960 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 886.050 3466.000 886.330 3470.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 4.000 786.720 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3451.720 4.000 3452.320 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 703.890 3466.000 704.170 3470.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2059.970 3466.000 2060.250 3470.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1663.450 3466.000 1663.730 3470.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.010 3466.000 323.290 3470.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1738.890 0.000 1739.170 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1574.210 0.000 1574.490 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3060.040 4.000 3060.640 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2106.680 4.000 2107.280 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1815.640 2700.000 1816.240 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 3457.360 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 3457.360 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.800 2694.220 3457.200 ;
      LAYER met1 ;
        RECT 5.520 4.460 2694.220 3457.360 ;
      LAYER met2 ;
        RECT 8.830 3465.720 9.010 3466.000 ;
        RECT 9.850 3465.720 25.570 3466.000 ;
        RECT 26.410 3465.720 42.130 3466.000 ;
        RECT 42.970 3465.720 58.690 3466.000 ;
        RECT 59.530 3465.720 75.250 3466.000 ;
        RECT 76.090 3465.720 91.810 3466.000 ;
        RECT 92.650 3465.720 108.370 3466.000 ;
        RECT 109.210 3465.720 124.930 3466.000 ;
        RECT 125.770 3465.720 141.490 3466.000 ;
        RECT 142.330 3465.720 158.050 3466.000 ;
        RECT 158.890 3465.720 174.610 3466.000 ;
        RECT 175.450 3465.720 190.250 3466.000 ;
        RECT 191.090 3465.720 206.810 3466.000 ;
        RECT 207.650 3465.720 223.370 3466.000 ;
        RECT 224.210 3465.720 239.930 3466.000 ;
        RECT 240.770 3465.720 256.490 3466.000 ;
        RECT 257.330 3465.720 273.050 3466.000 ;
        RECT 273.890 3465.720 289.610 3466.000 ;
        RECT 290.450 3465.720 306.170 3466.000 ;
        RECT 307.010 3465.720 322.730 3466.000 ;
        RECT 323.570 3465.720 339.290 3466.000 ;
        RECT 340.130 3465.720 355.850 3466.000 ;
        RECT 356.690 3465.720 372.410 3466.000 ;
        RECT 373.250 3465.720 388.970 3466.000 ;
        RECT 389.810 3465.720 405.530 3466.000 ;
        RECT 406.370 3465.720 422.090 3466.000 ;
        RECT 422.930 3465.720 438.650 3466.000 ;
        RECT 439.490 3465.720 455.210 3466.000 ;
        RECT 456.050 3465.720 471.770 3466.000 ;
        RECT 472.610 3465.720 488.330 3466.000 ;
        RECT 489.170 3465.720 504.890 3466.000 ;
        RECT 505.730 3465.720 521.450 3466.000 ;
        RECT 522.290 3465.720 538.010 3466.000 ;
        RECT 538.850 3465.720 554.570 3466.000 ;
        RECT 555.410 3465.720 571.130 3466.000 ;
        RECT 571.970 3465.720 587.690 3466.000 ;
        RECT 588.530 3465.720 604.250 3466.000 ;
        RECT 605.090 3465.720 620.810 3466.000 ;
        RECT 621.650 3465.720 637.370 3466.000 ;
        RECT 638.210 3465.720 653.930 3466.000 ;
        RECT 654.770 3465.720 670.490 3466.000 ;
        RECT 671.330 3465.720 687.050 3466.000 ;
        RECT 687.890 3465.720 703.610 3466.000 ;
        RECT 704.450 3465.720 720.170 3466.000 ;
        RECT 721.010 3465.720 736.730 3466.000 ;
        RECT 737.570 3465.720 753.290 3466.000 ;
        RECT 754.130 3465.720 769.850 3466.000 ;
        RECT 770.690 3465.720 786.410 3466.000 ;
        RECT 787.250 3465.720 802.970 3466.000 ;
        RECT 803.810 3465.720 819.530 3466.000 ;
        RECT 820.370 3465.720 836.090 3466.000 ;
        RECT 836.930 3465.720 852.650 3466.000 ;
        RECT 853.490 3465.720 869.210 3466.000 ;
        RECT 870.050 3465.720 885.770 3466.000 ;
        RECT 886.610 3465.720 902.330 3466.000 ;
        RECT 903.170 3465.720 918.890 3466.000 ;
        RECT 919.730 3465.720 935.450 3466.000 ;
        RECT 936.290 3465.720 952.010 3466.000 ;
        RECT 952.850 3465.720 968.570 3466.000 ;
        RECT 969.410 3465.720 985.130 3466.000 ;
        RECT 985.970 3465.720 1001.690 3466.000 ;
        RECT 1002.530 3465.720 1017.330 3466.000 ;
        RECT 1018.170 3465.720 1033.890 3466.000 ;
        RECT 1034.730 3465.720 1050.450 3466.000 ;
        RECT 1051.290 3465.720 1067.010 3466.000 ;
        RECT 1067.850 3465.720 1083.570 3466.000 ;
        RECT 1084.410 3465.720 1100.130 3466.000 ;
        RECT 1100.970 3465.720 1116.690 3466.000 ;
        RECT 1117.530 3465.720 1133.250 3466.000 ;
        RECT 1134.090 3465.720 1149.810 3466.000 ;
        RECT 1150.650 3465.720 1166.370 3466.000 ;
        RECT 1167.210 3465.720 1182.930 3466.000 ;
        RECT 1183.770 3465.720 1199.490 3466.000 ;
        RECT 1200.330 3465.720 1216.050 3466.000 ;
        RECT 1216.890 3465.720 1232.610 3466.000 ;
        RECT 1233.450 3465.720 1249.170 3466.000 ;
        RECT 1250.010 3465.720 1265.730 3466.000 ;
        RECT 1266.570 3465.720 1282.290 3466.000 ;
        RECT 1283.130 3465.720 1298.850 3466.000 ;
        RECT 1299.690 3465.720 1315.410 3466.000 ;
        RECT 1316.250 3465.720 1331.970 3466.000 ;
        RECT 1332.810 3465.720 1348.530 3466.000 ;
        RECT 1349.370 3465.720 1365.090 3466.000 ;
        RECT 1365.930 3465.720 1381.650 3466.000 ;
        RECT 1382.490 3465.720 1398.210 3466.000 ;
        RECT 1399.050 3465.720 1414.770 3466.000 ;
        RECT 1415.610 3465.720 1431.330 3466.000 ;
        RECT 1432.170 3465.720 1447.890 3466.000 ;
        RECT 1448.730 3465.720 1464.450 3466.000 ;
        RECT 1465.290 3465.720 1481.010 3466.000 ;
        RECT 1481.850 3465.720 1497.570 3466.000 ;
        RECT 1498.410 3465.720 1514.130 3466.000 ;
        RECT 1514.970 3465.720 1530.690 3466.000 ;
        RECT 1531.530 3465.720 1547.250 3466.000 ;
        RECT 1548.090 3465.720 1563.810 3466.000 ;
        RECT 1564.650 3465.720 1580.370 3466.000 ;
        RECT 1581.210 3465.720 1596.930 3466.000 ;
        RECT 1597.770 3465.720 1613.490 3466.000 ;
        RECT 1614.330 3465.720 1630.050 3466.000 ;
        RECT 1630.890 3465.720 1646.610 3466.000 ;
        RECT 1647.450 3465.720 1663.170 3466.000 ;
        RECT 1664.010 3465.720 1679.730 3466.000 ;
        RECT 1680.570 3465.720 1696.290 3466.000 ;
        RECT 1697.130 3465.720 1712.850 3466.000 ;
        RECT 1713.690 3465.720 1729.410 3466.000 ;
        RECT 1730.250 3465.720 1745.970 3466.000 ;
        RECT 1746.810 3465.720 1762.530 3466.000 ;
        RECT 1763.370 3465.720 1779.090 3466.000 ;
        RECT 1779.930 3465.720 1795.650 3466.000 ;
        RECT 1796.490 3465.720 1812.210 3466.000 ;
        RECT 1813.050 3465.720 1828.770 3466.000 ;
        RECT 1829.610 3465.720 1845.330 3466.000 ;
        RECT 1846.170 3465.720 1860.970 3466.000 ;
        RECT 1861.810 3465.720 1877.530 3466.000 ;
        RECT 1878.370 3465.720 1894.090 3466.000 ;
        RECT 1894.930 3465.720 1910.650 3466.000 ;
        RECT 1911.490 3465.720 1927.210 3466.000 ;
        RECT 1928.050 3465.720 1943.770 3466.000 ;
        RECT 1944.610 3465.720 1960.330 3466.000 ;
        RECT 1961.170 3465.720 1976.890 3466.000 ;
        RECT 1977.730 3465.720 1993.450 3466.000 ;
        RECT 1994.290 3465.720 2010.010 3466.000 ;
        RECT 2010.850 3465.720 2026.570 3466.000 ;
        RECT 2027.410 3465.720 2043.130 3466.000 ;
        RECT 2043.970 3465.720 2059.690 3466.000 ;
        RECT 2060.530 3465.720 2076.250 3466.000 ;
        RECT 2077.090 3465.720 2092.810 3466.000 ;
        RECT 2093.650 3465.720 2109.370 3466.000 ;
        RECT 2110.210 3465.720 2125.930 3466.000 ;
        RECT 2126.770 3465.720 2142.490 3466.000 ;
        RECT 2143.330 3465.720 2159.050 3466.000 ;
        RECT 2159.890 3465.720 2175.610 3466.000 ;
        RECT 2176.450 3465.720 2192.170 3466.000 ;
        RECT 2193.010 3465.720 2208.730 3466.000 ;
        RECT 2209.570 3465.720 2225.290 3466.000 ;
        RECT 2226.130 3465.720 2241.850 3466.000 ;
        RECT 2242.690 3465.720 2258.410 3466.000 ;
        RECT 2259.250 3465.720 2274.970 3466.000 ;
        RECT 2275.810 3465.720 2291.530 3466.000 ;
        RECT 2292.370 3465.720 2308.090 3466.000 ;
        RECT 2308.930 3465.720 2324.650 3466.000 ;
        RECT 2325.490 3465.720 2341.210 3466.000 ;
        RECT 2342.050 3465.720 2357.770 3466.000 ;
        RECT 2358.610 3465.720 2374.330 3466.000 ;
        RECT 2375.170 3465.720 2390.890 3466.000 ;
        RECT 2391.730 3465.720 2407.450 3466.000 ;
        RECT 2408.290 3465.720 2424.010 3466.000 ;
        RECT 2424.850 3465.720 2440.570 3466.000 ;
        RECT 2441.410 3465.720 2457.130 3466.000 ;
        RECT 2457.970 3465.720 2473.690 3466.000 ;
        RECT 2474.530 3465.720 2490.250 3466.000 ;
        RECT 2491.090 3465.720 2506.810 3466.000 ;
        RECT 2507.650 3465.720 2523.370 3466.000 ;
        RECT 2524.210 3465.720 2539.930 3466.000 ;
        RECT 2540.770 3465.720 2556.490 3466.000 ;
        RECT 2557.330 3465.720 2573.050 3466.000 ;
        RECT 2573.890 3465.720 2589.610 3466.000 ;
        RECT 2590.450 3465.720 2606.170 3466.000 ;
        RECT 2607.010 3465.720 2622.730 3466.000 ;
        RECT 2623.570 3465.720 2639.290 3466.000 ;
        RECT 2640.130 3465.720 2655.850 3466.000 ;
        RECT 2656.690 3465.720 2672.410 3466.000 ;
        RECT 2673.250 3465.720 2687.690 3466.000 ;
        RECT 8.830 4.280 2687.690 3465.720 ;
        RECT 8.830 4.000 18.210 4.280 ;
        RECT 19.050 4.000 34.770 4.280 ;
        RECT 35.610 4.000 51.330 4.280 ;
        RECT 52.170 4.000 67.890 4.280 ;
        RECT 68.730 4.000 84.450 4.280 ;
        RECT 85.290 4.000 101.010 4.280 ;
        RECT 101.850 4.000 117.570 4.280 ;
        RECT 118.410 4.000 134.130 4.280 ;
        RECT 134.970 4.000 150.690 4.280 ;
        RECT 151.530 4.000 167.250 4.280 ;
        RECT 168.090 4.000 183.810 4.280 ;
        RECT 184.650 4.000 200.370 4.280 ;
        RECT 201.210 4.000 216.930 4.280 ;
        RECT 217.770 4.000 233.490 4.280 ;
        RECT 234.330 4.000 250.050 4.280 ;
        RECT 250.890 4.000 266.610 4.280 ;
        RECT 267.450 4.000 283.170 4.280 ;
        RECT 284.010 4.000 299.730 4.280 ;
        RECT 300.570 4.000 316.290 4.280 ;
        RECT 317.130 4.000 332.850 4.280 ;
        RECT 333.690 4.000 349.410 4.280 ;
        RECT 350.250 4.000 365.970 4.280 ;
        RECT 366.810 4.000 382.530 4.280 ;
        RECT 383.370 4.000 399.090 4.280 ;
        RECT 399.930 4.000 415.650 4.280 ;
        RECT 416.490 4.000 432.210 4.280 ;
        RECT 433.050 4.000 448.770 4.280 ;
        RECT 449.610 4.000 465.330 4.280 ;
        RECT 466.170 4.000 481.890 4.280 ;
        RECT 482.730 4.000 498.450 4.280 ;
        RECT 499.290 4.000 515.010 4.280 ;
        RECT 515.850 4.000 531.570 4.280 ;
        RECT 532.410 4.000 548.130 4.280 ;
        RECT 548.970 4.000 564.690 4.280 ;
        RECT 565.530 4.000 581.250 4.280 ;
        RECT 582.090 4.000 597.810 4.280 ;
        RECT 598.650 4.000 614.370 4.280 ;
        RECT 615.210 4.000 630.930 4.280 ;
        RECT 631.770 4.000 647.490 4.280 ;
        RECT 648.330 4.000 664.050 4.280 ;
        RECT 664.890 4.000 680.610 4.280 ;
        RECT 681.450 4.000 697.170 4.280 ;
        RECT 698.010 4.000 713.730 4.280 ;
        RECT 714.570 4.000 730.290 4.280 ;
        RECT 731.130 4.000 746.850 4.280 ;
        RECT 747.690 4.000 763.410 4.280 ;
        RECT 764.250 4.000 779.970 4.280 ;
        RECT 780.810 4.000 796.530 4.280 ;
        RECT 797.370 4.000 813.090 4.280 ;
        RECT 813.930 4.000 829.650 4.280 ;
        RECT 830.490 4.000 845.290 4.280 ;
        RECT 846.130 4.000 861.850 4.280 ;
        RECT 862.690 4.000 878.410 4.280 ;
        RECT 879.250 4.000 894.970 4.280 ;
        RECT 895.810 4.000 911.530 4.280 ;
        RECT 912.370 4.000 928.090 4.280 ;
        RECT 928.930 4.000 944.650 4.280 ;
        RECT 945.490 4.000 961.210 4.280 ;
        RECT 962.050 4.000 977.770 4.280 ;
        RECT 978.610 4.000 994.330 4.280 ;
        RECT 995.170 4.000 1010.890 4.280 ;
        RECT 1011.730 4.000 1027.450 4.280 ;
        RECT 1028.290 4.000 1044.010 4.280 ;
        RECT 1044.850 4.000 1060.570 4.280 ;
        RECT 1061.410 4.000 1077.130 4.280 ;
        RECT 1077.970 4.000 1093.690 4.280 ;
        RECT 1094.530 4.000 1110.250 4.280 ;
        RECT 1111.090 4.000 1126.810 4.280 ;
        RECT 1127.650 4.000 1143.370 4.280 ;
        RECT 1144.210 4.000 1159.930 4.280 ;
        RECT 1160.770 4.000 1176.490 4.280 ;
        RECT 1177.330 4.000 1193.050 4.280 ;
        RECT 1193.890 4.000 1209.610 4.280 ;
        RECT 1210.450 4.000 1226.170 4.280 ;
        RECT 1227.010 4.000 1242.730 4.280 ;
        RECT 1243.570 4.000 1259.290 4.280 ;
        RECT 1260.130 4.000 1275.850 4.280 ;
        RECT 1276.690 4.000 1292.410 4.280 ;
        RECT 1293.250 4.000 1308.970 4.280 ;
        RECT 1309.810 4.000 1325.530 4.280 ;
        RECT 1326.370 4.000 1342.090 4.280 ;
        RECT 1342.930 4.000 1358.650 4.280 ;
        RECT 1359.490 4.000 1375.210 4.280 ;
        RECT 1376.050 4.000 1391.770 4.280 ;
        RECT 1392.610 4.000 1408.330 4.280 ;
        RECT 1409.170 4.000 1424.890 4.280 ;
        RECT 1425.730 4.000 1441.450 4.280 ;
        RECT 1442.290 4.000 1458.010 4.280 ;
        RECT 1458.850 4.000 1474.570 4.280 ;
        RECT 1475.410 4.000 1491.130 4.280 ;
        RECT 1491.970 4.000 1507.690 4.280 ;
        RECT 1508.530 4.000 1524.250 4.280 ;
        RECT 1525.090 4.000 1540.810 4.280 ;
        RECT 1541.650 4.000 1557.370 4.280 ;
        RECT 1558.210 4.000 1573.930 4.280 ;
        RECT 1574.770 4.000 1590.490 4.280 ;
        RECT 1591.330 4.000 1607.050 4.280 ;
        RECT 1607.890 4.000 1623.610 4.280 ;
        RECT 1624.450 4.000 1640.170 4.280 ;
        RECT 1641.010 4.000 1656.730 4.280 ;
        RECT 1657.570 4.000 1673.290 4.280 ;
        RECT 1674.130 4.000 1688.930 4.280 ;
        RECT 1689.770 4.000 1705.490 4.280 ;
        RECT 1706.330 4.000 1722.050 4.280 ;
        RECT 1722.890 4.000 1738.610 4.280 ;
        RECT 1739.450 4.000 1755.170 4.280 ;
        RECT 1756.010 4.000 1771.730 4.280 ;
        RECT 1772.570 4.000 1788.290 4.280 ;
        RECT 1789.130 4.000 1804.850 4.280 ;
        RECT 1805.690 4.000 1821.410 4.280 ;
        RECT 1822.250 4.000 1837.970 4.280 ;
        RECT 1838.810 4.000 1854.530 4.280 ;
        RECT 1855.370 4.000 1871.090 4.280 ;
        RECT 1871.930 4.000 1887.650 4.280 ;
        RECT 1888.490 4.000 1904.210 4.280 ;
        RECT 1905.050 4.000 1920.770 4.280 ;
        RECT 1921.610 4.000 1937.330 4.280 ;
        RECT 1938.170 4.000 1953.890 4.280 ;
        RECT 1954.730 4.000 1970.450 4.280 ;
        RECT 1971.290 4.000 1987.010 4.280 ;
        RECT 1987.850 4.000 2003.570 4.280 ;
        RECT 2004.410 4.000 2020.130 4.280 ;
        RECT 2020.970 4.000 2036.690 4.280 ;
        RECT 2037.530 4.000 2053.250 4.280 ;
        RECT 2054.090 4.000 2069.810 4.280 ;
        RECT 2070.650 4.000 2086.370 4.280 ;
        RECT 2087.210 4.000 2102.930 4.280 ;
        RECT 2103.770 4.000 2119.490 4.280 ;
        RECT 2120.330 4.000 2136.050 4.280 ;
        RECT 2136.890 4.000 2152.610 4.280 ;
        RECT 2153.450 4.000 2169.170 4.280 ;
        RECT 2170.010 4.000 2185.730 4.280 ;
        RECT 2186.570 4.000 2202.290 4.280 ;
        RECT 2203.130 4.000 2218.850 4.280 ;
        RECT 2219.690 4.000 2235.410 4.280 ;
        RECT 2236.250 4.000 2251.970 4.280 ;
        RECT 2252.810 4.000 2268.530 4.280 ;
        RECT 2269.370 4.000 2285.090 4.280 ;
        RECT 2285.930 4.000 2301.650 4.280 ;
        RECT 2302.490 4.000 2318.210 4.280 ;
        RECT 2319.050 4.000 2334.770 4.280 ;
        RECT 2335.610 4.000 2351.330 4.280 ;
        RECT 2352.170 4.000 2367.890 4.280 ;
        RECT 2368.730 4.000 2384.450 4.280 ;
        RECT 2385.290 4.000 2401.010 4.280 ;
        RECT 2401.850 4.000 2417.570 4.280 ;
        RECT 2418.410 4.000 2434.130 4.280 ;
        RECT 2434.970 4.000 2450.690 4.280 ;
        RECT 2451.530 4.000 2467.250 4.280 ;
        RECT 2468.090 4.000 2483.810 4.280 ;
        RECT 2484.650 4.000 2500.370 4.280 ;
        RECT 2501.210 4.000 2516.930 4.280 ;
        RECT 2517.770 4.000 2532.570 4.280 ;
        RECT 2533.410 4.000 2549.130 4.280 ;
        RECT 2549.970 4.000 2565.690 4.280 ;
        RECT 2566.530 4.000 2582.250 4.280 ;
        RECT 2583.090 4.000 2598.810 4.280 ;
        RECT 2599.650 4.000 2615.370 4.280 ;
        RECT 2616.210 4.000 2631.930 4.280 ;
        RECT 2632.770 4.000 2648.490 4.280 ;
        RECT 2649.330 4.000 2665.050 4.280 ;
        RECT 2665.890 4.000 2681.610 4.280 ;
        RECT 2682.450 4.000 2687.690 4.280 ;
      LAYER met3 ;
        RECT 3.990 3455.440 2696.000 3457.285 ;
        RECT 3.990 3454.040 2695.600 3455.440 ;
        RECT 3.990 3452.720 2696.000 3454.040 ;
        RECT 4.400 3451.320 2696.000 3452.720 ;
        RECT 3.990 3430.960 2696.000 3451.320 ;
        RECT 3.990 3429.560 2695.600 3430.960 ;
        RECT 3.990 3428.240 2696.000 3429.560 ;
        RECT 4.400 3426.840 2696.000 3428.240 ;
        RECT 3.990 3406.480 2696.000 3426.840 ;
        RECT 3.990 3405.080 2695.600 3406.480 ;
        RECT 3.990 3403.760 2696.000 3405.080 ;
        RECT 4.400 3402.360 2696.000 3403.760 ;
        RECT 3.990 3382.000 2696.000 3402.360 ;
        RECT 3.990 3380.600 2695.600 3382.000 ;
        RECT 3.990 3379.280 2696.000 3380.600 ;
        RECT 4.400 3377.880 2696.000 3379.280 ;
        RECT 3.990 3357.520 2696.000 3377.880 ;
        RECT 3.990 3356.120 2695.600 3357.520 ;
        RECT 3.990 3354.800 2696.000 3356.120 ;
        RECT 4.400 3353.400 2696.000 3354.800 ;
        RECT 3.990 3333.040 2696.000 3353.400 ;
        RECT 3.990 3331.640 2695.600 3333.040 ;
        RECT 3.990 3330.320 2696.000 3331.640 ;
        RECT 4.400 3328.920 2696.000 3330.320 ;
        RECT 3.990 3308.560 2696.000 3328.920 ;
        RECT 3.990 3307.160 2695.600 3308.560 ;
        RECT 3.990 3305.840 2696.000 3307.160 ;
        RECT 4.400 3304.440 2696.000 3305.840 ;
        RECT 3.990 3284.080 2696.000 3304.440 ;
        RECT 3.990 3282.680 2695.600 3284.080 ;
        RECT 3.990 3281.360 2696.000 3282.680 ;
        RECT 4.400 3279.960 2696.000 3281.360 ;
        RECT 3.990 3259.600 2696.000 3279.960 ;
        RECT 3.990 3258.200 2695.600 3259.600 ;
        RECT 3.990 3256.880 2696.000 3258.200 ;
        RECT 4.400 3255.480 2696.000 3256.880 ;
        RECT 3.990 3235.120 2696.000 3255.480 ;
        RECT 3.990 3233.720 2695.600 3235.120 ;
        RECT 3.990 3232.400 2696.000 3233.720 ;
        RECT 4.400 3231.000 2696.000 3232.400 ;
        RECT 3.990 3210.640 2696.000 3231.000 ;
        RECT 3.990 3209.240 2695.600 3210.640 ;
        RECT 3.990 3207.920 2696.000 3209.240 ;
        RECT 4.400 3206.520 2696.000 3207.920 ;
        RECT 3.990 3186.160 2696.000 3206.520 ;
        RECT 3.990 3184.760 2695.600 3186.160 ;
        RECT 3.990 3183.440 2696.000 3184.760 ;
        RECT 4.400 3182.040 2696.000 3183.440 ;
        RECT 3.990 3161.680 2696.000 3182.040 ;
        RECT 3.990 3160.280 2695.600 3161.680 ;
        RECT 3.990 3158.960 2696.000 3160.280 ;
        RECT 4.400 3157.560 2696.000 3158.960 ;
        RECT 3.990 3137.200 2696.000 3157.560 ;
        RECT 3.990 3135.800 2695.600 3137.200 ;
        RECT 3.990 3134.480 2696.000 3135.800 ;
        RECT 4.400 3133.080 2696.000 3134.480 ;
        RECT 3.990 3112.720 2696.000 3133.080 ;
        RECT 3.990 3111.320 2695.600 3112.720 ;
        RECT 3.990 3110.000 2696.000 3111.320 ;
        RECT 4.400 3108.600 2696.000 3110.000 ;
        RECT 3.990 3088.240 2696.000 3108.600 ;
        RECT 3.990 3086.840 2695.600 3088.240 ;
        RECT 3.990 3085.520 2696.000 3086.840 ;
        RECT 4.400 3084.120 2696.000 3085.520 ;
        RECT 3.990 3063.760 2696.000 3084.120 ;
        RECT 3.990 3062.360 2695.600 3063.760 ;
        RECT 3.990 3061.040 2696.000 3062.360 ;
        RECT 4.400 3059.640 2696.000 3061.040 ;
        RECT 3.990 3039.280 2696.000 3059.640 ;
        RECT 3.990 3037.880 2695.600 3039.280 ;
        RECT 3.990 3036.560 2696.000 3037.880 ;
        RECT 4.400 3035.160 2696.000 3036.560 ;
        RECT 3.990 3014.800 2696.000 3035.160 ;
        RECT 3.990 3013.400 2695.600 3014.800 ;
        RECT 3.990 3012.080 2696.000 3013.400 ;
        RECT 4.400 3010.680 2696.000 3012.080 ;
        RECT 3.990 2990.320 2696.000 3010.680 ;
        RECT 3.990 2988.920 2695.600 2990.320 ;
        RECT 3.990 2987.600 2696.000 2988.920 ;
        RECT 4.400 2986.200 2696.000 2987.600 ;
        RECT 3.990 2965.840 2696.000 2986.200 ;
        RECT 3.990 2964.440 2695.600 2965.840 ;
        RECT 3.990 2963.120 2696.000 2964.440 ;
        RECT 4.400 2961.720 2696.000 2963.120 ;
        RECT 3.990 2941.360 2696.000 2961.720 ;
        RECT 3.990 2939.960 2695.600 2941.360 ;
        RECT 3.990 2938.640 2696.000 2939.960 ;
        RECT 4.400 2937.240 2696.000 2938.640 ;
        RECT 3.990 2916.880 2696.000 2937.240 ;
        RECT 3.990 2915.480 2695.600 2916.880 ;
        RECT 3.990 2914.160 2696.000 2915.480 ;
        RECT 4.400 2912.760 2696.000 2914.160 ;
        RECT 3.990 2892.400 2696.000 2912.760 ;
        RECT 3.990 2891.000 2695.600 2892.400 ;
        RECT 3.990 2889.680 2696.000 2891.000 ;
        RECT 4.400 2888.280 2696.000 2889.680 ;
        RECT 3.990 2867.920 2696.000 2888.280 ;
        RECT 3.990 2866.520 2695.600 2867.920 ;
        RECT 3.990 2865.200 2696.000 2866.520 ;
        RECT 4.400 2863.800 2696.000 2865.200 ;
        RECT 3.990 2843.440 2696.000 2863.800 ;
        RECT 3.990 2842.040 2695.600 2843.440 ;
        RECT 3.990 2840.720 2696.000 2842.040 ;
        RECT 4.400 2839.320 2696.000 2840.720 ;
        RECT 3.990 2818.960 2696.000 2839.320 ;
        RECT 3.990 2817.560 2695.600 2818.960 ;
        RECT 3.990 2816.240 2696.000 2817.560 ;
        RECT 4.400 2814.840 2696.000 2816.240 ;
        RECT 3.990 2794.480 2696.000 2814.840 ;
        RECT 3.990 2793.080 2695.600 2794.480 ;
        RECT 3.990 2791.760 2696.000 2793.080 ;
        RECT 4.400 2790.360 2696.000 2791.760 ;
        RECT 3.990 2770.000 2696.000 2790.360 ;
        RECT 3.990 2768.600 2695.600 2770.000 ;
        RECT 3.990 2767.280 2696.000 2768.600 ;
        RECT 4.400 2765.880 2696.000 2767.280 ;
        RECT 3.990 2745.520 2696.000 2765.880 ;
        RECT 3.990 2744.120 2695.600 2745.520 ;
        RECT 3.990 2742.800 2696.000 2744.120 ;
        RECT 4.400 2741.400 2696.000 2742.800 ;
        RECT 3.990 2721.040 2696.000 2741.400 ;
        RECT 3.990 2719.640 2695.600 2721.040 ;
        RECT 3.990 2718.320 2696.000 2719.640 ;
        RECT 4.400 2716.920 2696.000 2718.320 ;
        RECT 3.990 2696.560 2696.000 2716.920 ;
        RECT 3.990 2695.160 2695.600 2696.560 ;
        RECT 3.990 2693.840 2696.000 2695.160 ;
        RECT 4.400 2692.440 2696.000 2693.840 ;
        RECT 3.990 2672.080 2696.000 2692.440 ;
        RECT 3.990 2670.680 2695.600 2672.080 ;
        RECT 3.990 2669.360 2696.000 2670.680 ;
        RECT 4.400 2667.960 2696.000 2669.360 ;
        RECT 3.990 2647.600 2696.000 2667.960 ;
        RECT 3.990 2646.200 2695.600 2647.600 ;
        RECT 3.990 2644.880 2696.000 2646.200 ;
        RECT 4.400 2643.480 2696.000 2644.880 ;
        RECT 3.990 2623.120 2696.000 2643.480 ;
        RECT 3.990 2621.720 2695.600 2623.120 ;
        RECT 3.990 2620.400 2696.000 2621.720 ;
        RECT 4.400 2619.000 2696.000 2620.400 ;
        RECT 3.990 2598.640 2696.000 2619.000 ;
        RECT 3.990 2597.240 2695.600 2598.640 ;
        RECT 3.990 2595.920 2696.000 2597.240 ;
        RECT 4.400 2594.520 2696.000 2595.920 ;
        RECT 3.990 2574.160 2696.000 2594.520 ;
        RECT 3.990 2572.760 2695.600 2574.160 ;
        RECT 3.990 2571.440 2696.000 2572.760 ;
        RECT 4.400 2570.040 2696.000 2571.440 ;
        RECT 3.990 2549.680 2696.000 2570.040 ;
        RECT 3.990 2548.280 2695.600 2549.680 ;
        RECT 3.990 2546.960 2696.000 2548.280 ;
        RECT 4.400 2545.560 2696.000 2546.960 ;
        RECT 3.990 2525.200 2696.000 2545.560 ;
        RECT 3.990 2523.800 2695.600 2525.200 ;
        RECT 3.990 2522.480 2696.000 2523.800 ;
        RECT 4.400 2521.080 2696.000 2522.480 ;
        RECT 3.990 2500.720 2696.000 2521.080 ;
        RECT 3.990 2499.320 2695.600 2500.720 ;
        RECT 3.990 2498.000 2696.000 2499.320 ;
        RECT 4.400 2496.600 2696.000 2498.000 ;
        RECT 3.990 2476.240 2696.000 2496.600 ;
        RECT 3.990 2474.880 2695.600 2476.240 ;
        RECT 4.400 2474.840 2695.600 2474.880 ;
        RECT 4.400 2473.480 2696.000 2474.840 ;
        RECT 3.990 2451.760 2696.000 2473.480 ;
        RECT 3.990 2450.400 2695.600 2451.760 ;
        RECT 4.400 2450.360 2695.600 2450.400 ;
        RECT 4.400 2449.000 2696.000 2450.360 ;
        RECT 3.990 2427.280 2696.000 2449.000 ;
        RECT 3.990 2425.920 2695.600 2427.280 ;
        RECT 4.400 2425.880 2695.600 2425.920 ;
        RECT 4.400 2424.520 2696.000 2425.880 ;
        RECT 3.990 2402.800 2696.000 2424.520 ;
        RECT 3.990 2401.440 2695.600 2402.800 ;
        RECT 4.400 2401.400 2695.600 2401.440 ;
        RECT 4.400 2400.040 2696.000 2401.400 ;
        RECT 3.990 2378.320 2696.000 2400.040 ;
        RECT 3.990 2376.960 2695.600 2378.320 ;
        RECT 4.400 2376.920 2695.600 2376.960 ;
        RECT 4.400 2375.560 2696.000 2376.920 ;
        RECT 3.990 2353.840 2696.000 2375.560 ;
        RECT 3.990 2352.480 2695.600 2353.840 ;
        RECT 4.400 2352.440 2695.600 2352.480 ;
        RECT 4.400 2351.080 2696.000 2352.440 ;
        RECT 3.990 2329.360 2696.000 2351.080 ;
        RECT 3.990 2328.000 2695.600 2329.360 ;
        RECT 4.400 2327.960 2695.600 2328.000 ;
        RECT 4.400 2326.600 2696.000 2327.960 ;
        RECT 3.990 2304.880 2696.000 2326.600 ;
        RECT 3.990 2303.520 2695.600 2304.880 ;
        RECT 4.400 2303.480 2695.600 2303.520 ;
        RECT 4.400 2302.120 2696.000 2303.480 ;
        RECT 3.990 2280.400 2696.000 2302.120 ;
        RECT 3.990 2279.040 2695.600 2280.400 ;
        RECT 4.400 2279.000 2695.600 2279.040 ;
        RECT 4.400 2277.640 2696.000 2279.000 ;
        RECT 3.990 2255.920 2696.000 2277.640 ;
        RECT 3.990 2254.560 2695.600 2255.920 ;
        RECT 4.400 2254.520 2695.600 2254.560 ;
        RECT 4.400 2253.160 2696.000 2254.520 ;
        RECT 3.990 2231.440 2696.000 2253.160 ;
        RECT 3.990 2230.080 2695.600 2231.440 ;
        RECT 4.400 2230.040 2695.600 2230.080 ;
        RECT 4.400 2228.680 2696.000 2230.040 ;
        RECT 3.990 2208.320 2696.000 2228.680 ;
        RECT 3.990 2206.920 2695.600 2208.320 ;
        RECT 3.990 2205.600 2696.000 2206.920 ;
        RECT 4.400 2204.200 2696.000 2205.600 ;
        RECT 3.990 2183.840 2696.000 2204.200 ;
        RECT 3.990 2182.440 2695.600 2183.840 ;
        RECT 3.990 2181.120 2696.000 2182.440 ;
        RECT 4.400 2179.720 2696.000 2181.120 ;
        RECT 3.990 2159.360 2696.000 2179.720 ;
        RECT 3.990 2157.960 2695.600 2159.360 ;
        RECT 3.990 2156.640 2696.000 2157.960 ;
        RECT 4.400 2155.240 2696.000 2156.640 ;
        RECT 3.990 2134.880 2696.000 2155.240 ;
        RECT 3.990 2133.480 2695.600 2134.880 ;
        RECT 3.990 2132.160 2696.000 2133.480 ;
        RECT 4.400 2130.760 2696.000 2132.160 ;
        RECT 3.990 2110.400 2696.000 2130.760 ;
        RECT 3.990 2109.000 2695.600 2110.400 ;
        RECT 3.990 2107.680 2696.000 2109.000 ;
        RECT 4.400 2106.280 2696.000 2107.680 ;
        RECT 3.990 2085.920 2696.000 2106.280 ;
        RECT 3.990 2084.520 2695.600 2085.920 ;
        RECT 3.990 2083.200 2696.000 2084.520 ;
        RECT 4.400 2081.800 2696.000 2083.200 ;
        RECT 3.990 2061.440 2696.000 2081.800 ;
        RECT 3.990 2060.040 2695.600 2061.440 ;
        RECT 3.990 2058.720 2696.000 2060.040 ;
        RECT 4.400 2057.320 2696.000 2058.720 ;
        RECT 3.990 2036.960 2696.000 2057.320 ;
        RECT 3.990 2035.560 2695.600 2036.960 ;
        RECT 3.990 2034.240 2696.000 2035.560 ;
        RECT 4.400 2032.840 2696.000 2034.240 ;
        RECT 3.990 2012.480 2696.000 2032.840 ;
        RECT 3.990 2011.080 2695.600 2012.480 ;
        RECT 3.990 2009.760 2696.000 2011.080 ;
        RECT 4.400 2008.360 2696.000 2009.760 ;
        RECT 3.990 1988.000 2696.000 2008.360 ;
        RECT 3.990 1986.600 2695.600 1988.000 ;
        RECT 3.990 1985.280 2696.000 1986.600 ;
        RECT 4.400 1983.880 2696.000 1985.280 ;
        RECT 3.990 1963.520 2696.000 1983.880 ;
        RECT 3.990 1962.120 2695.600 1963.520 ;
        RECT 3.990 1960.800 2696.000 1962.120 ;
        RECT 4.400 1959.400 2696.000 1960.800 ;
        RECT 3.990 1939.040 2696.000 1959.400 ;
        RECT 3.990 1937.640 2695.600 1939.040 ;
        RECT 3.990 1936.320 2696.000 1937.640 ;
        RECT 4.400 1934.920 2696.000 1936.320 ;
        RECT 3.990 1914.560 2696.000 1934.920 ;
        RECT 3.990 1913.160 2695.600 1914.560 ;
        RECT 3.990 1911.840 2696.000 1913.160 ;
        RECT 4.400 1910.440 2696.000 1911.840 ;
        RECT 3.990 1890.080 2696.000 1910.440 ;
        RECT 3.990 1888.680 2695.600 1890.080 ;
        RECT 3.990 1887.360 2696.000 1888.680 ;
        RECT 4.400 1885.960 2696.000 1887.360 ;
        RECT 3.990 1865.600 2696.000 1885.960 ;
        RECT 3.990 1864.200 2695.600 1865.600 ;
        RECT 3.990 1862.880 2696.000 1864.200 ;
        RECT 4.400 1861.480 2696.000 1862.880 ;
        RECT 3.990 1841.120 2696.000 1861.480 ;
        RECT 3.990 1839.720 2695.600 1841.120 ;
        RECT 3.990 1838.400 2696.000 1839.720 ;
        RECT 4.400 1837.000 2696.000 1838.400 ;
        RECT 3.990 1816.640 2696.000 1837.000 ;
        RECT 3.990 1815.240 2695.600 1816.640 ;
        RECT 3.990 1813.920 2696.000 1815.240 ;
        RECT 4.400 1812.520 2696.000 1813.920 ;
        RECT 3.990 1792.160 2696.000 1812.520 ;
        RECT 3.990 1790.760 2695.600 1792.160 ;
        RECT 3.990 1789.440 2696.000 1790.760 ;
        RECT 4.400 1788.040 2696.000 1789.440 ;
        RECT 3.990 1767.680 2696.000 1788.040 ;
        RECT 3.990 1766.280 2695.600 1767.680 ;
        RECT 3.990 1764.960 2696.000 1766.280 ;
        RECT 4.400 1763.560 2696.000 1764.960 ;
        RECT 3.990 1743.200 2696.000 1763.560 ;
        RECT 3.990 1741.800 2695.600 1743.200 ;
        RECT 3.990 1740.480 2696.000 1741.800 ;
        RECT 4.400 1739.080 2696.000 1740.480 ;
        RECT 3.990 1718.720 2696.000 1739.080 ;
        RECT 3.990 1717.320 2695.600 1718.720 ;
        RECT 3.990 1716.000 2696.000 1717.320 ;
        RECT 4.400 1714.600 2696.000 1716.000 ;
        RECT 3.990 1694.240 2696.000 1714.600 ;
        RECT 3.990 1692.840 2695.600 1694.240 ;
        RECT 3.990 1691.520 2696.000 1692.840 ;
        RECT 4.400 1690.120 2696.000 1691.520 ;
        RECT 3.990 1669.760 2696.000 1690.120 ;
        RECT 3.990 1668.360 2695.600 1669.760 ;
        RECT 3.990 1667.040 2696.000 1668.360 ;
        RECT 4.400 1665.640 2696.000 1667.040 ;
        RECT 3.990 1645.280 2696.000 1665.640 ;
        RECT 3.990 1643.880 2695.600 1645.280 ;
        RECT 3.990 1642.560 2696.000 1643.880 ;
        RECT 4.400 1641.160 2696.000 1642.560 ;
        RECT 3.990 1620.800 2696.000 1641.160 ;
        RECT 3.990 1619.400 2695.600 1620.800 ;
        RECT 3.990 1618.080 2696.000 1619.400 ;
        RECT 4.400 1616.680 2696.000 1618.080 ;
        RECT 3.990 1596.320 2696.000 1616.680 ;
        RECT 3.990 1594.920 2695.600 1596.320 ;
        RECT 3.990 1593.600 2696.000 1594.920 ;
        RECT 4.400 1592.200 2696.000 1593.600 ;
        RECT 3.990 1571.840 2696.000 1592.200 ;
        RECT 3.990 1570.440 2695.600 1571.840 ;
        RECT 3.990 1569.120 2696.000 1570.440 ;
        RECT 4.400 1567.720 2696.000 1569.120 ;
        RECT 3.990 1547.360 2696.000 1567.720 ;
        RECT 3.990 1545.960 2695.600 1547.360 ;
        RECT 3.990 1544.640 2696.000 1545.960 ;
        RECT 4.400 1543.240 2696.000 1544.640 ;
        RECT 3.990 1522.880 2696.000 1543.240 ;
        RECT 3.990 1521.480 2695.600 1522.880 ;
        RECT 3.990 1520.160 2696.000 1521.480 ;
        RECT 4.400 1518.760 2696.000 1520.160 ;
        RECT 3.990 1498.400 2696.000 1518.760 ;
        RECT 3.990 1497.000 2695.600 1498.400 ;
        RECT 3.990 1495.680 2696.000 1497.000 ;
        RECT 4.400 1494.280 2696.000 1495.680 ;
        RECT 3.990 1473.920 2696.000 1494.280 ;
        RECT 3.990 1472.520 2695.600 1473.920 ;
        RECT 3.990 1471.200 2696.000 1472.520 ;
        RECT 4.400 1469.800 2696.000 1471.200 ;
        RECT 3.990 1449.440 2696.000 1469.800 ;
        RECT 3.990 1448.040 2695.600 1449.440 ;
        RECT 3.990 1446.720 2696.000 1448.040 ;
        RECT 4.400 1445.320 2696.000 1446.720 ;
        RECT 3.990 1424.960 2696.000 1445.320 ;
        RECT 3.990 1423.560 2695.600 1424.960 ;
        RECT 3.990 1422.240 2696.000 1423.560 ;
        RECT 4.400 1420.840 2696.000 1422.240 ;
        RECT 3.990 1400.480 2696.000 1420.840 ;
        RECT 3.990 1399.080 2695.600 1400.480 ;
        RECT 3.990 1397.760 2696.000 1399.080 ;
        RECT 4.400 1396.360 2696.000 1397.760 ;
        RECT 3.990 1376.000 2696.000 1396.360 ;
        RECT 3.990 1374.600 2695.600 1376.000 ;
        RECT 3.990 1373.280 2696.000 1374.600 ;
        RECT 4.400 1371.880 2696.000 1373.280 ;
        RECT 3.990 1351.520 2696.000 1371.880 ;
        RECT 3.990 1350.120 2695.600 1351.520 ;
        RECT 3.990 1348.800 2696.000 1350.120 ;
        RECT 4.400 1347.400 2696.000 1348.800 ;
        RECT 3.990 1327.040 2696.000 1347.400 ;
        RECT 3.990 1325.640 2695.600 1327.040 ;
        RECT 3.990 1324.320 2696.000 1325.640 ;
        RECT 4.400 1322.920 2696.000 1324.320 ;
        RECT 3.990 1302.560 2696.000 1322.920 ;
        RECT 3.990 1301.160 2695.600 1302.560 ;
        RECT 3.990 1299.840 2696.000 1301.160 ;
        RECT 4.400 1298.440 2696.000 1299.840 ;
        RECT 3.990 1278.080 2696.000 1298.440 ;
        RECT 3.990 1276.680 2695.600 1278.080 ;
        RECT 3.990 1275.360 2696.000 1276.680 ;
        RECT 4.400 1273.960 2696.000 1275.360 ;
        RECT 3.990 1253.600 2696.000 1273.960 ;
        RECT 3.990 1252.200 2695.600 1253.600 ;
        RECT 3.990 1250.880 2696.000 1252.200 ;
        RECT 4.400 1249.480 2696.000 1250.880 ;
        RECT 3.990 1229.120 2696.000 1249.480 ;
        RECT 3.990 1227.760 2695.600 1229.120 ;
        RECT 4.400 1227.720 2695.600 1227.760 ;
        RECT 4.400 1226.360 2696.000 1227.720 ;
        RECT 3.990 1204.640 2696.000 1226.360 ;
        RECT 3.990 1203.280 2695.600 1204.640 ;
        RECT 4.400 1203.240 2695.600 1203.280 ;
        RECT 4.400 1201.880 2696.000 1203.240 ;
        RECT 3.990 1180.160 2696.000 1201.880 ;
        RECT 3.990 1178.800 2695.600 1180.160 ;
        RECT 4.400 1178.760 2695.600 1178.800 ;
        RECT 4.400 1177.400 2696.000 1178.760 ;
        RECT 3.990 1155.680 2696.000 1177.400 ;
        RECT 3.990 1154.320 2695.600 1155.680 ;
        RECT 4.400 1154.280 2695.600 1154.320 ;
        RECT 4.400 1152.920 2696.000 1154.280 ;
        RECT 3.990 1131.200 2696.000 1152.920 ;
        RECT 3.990 1129.840 2695.600 1131.200 ;
        RECT 4.400 1129.800 2695.600 1129.840 ;
        RECT 4.400 1128.440 2696.000 1129.800 ;
        RECT 3.990 1106.720 2696.000 1128.440 ;
        RECT 3.990 1105.360 2695.600 1106.720 ;
        RECT 4.400 1105.320 2695.600 1105.360 ;
        RECT 4.400 1103.960 2696.000 1105.320 ;
        RECT 3.990 1082.240 2696.000 1103.960 ;
        RECT 3.990 1080.880 2695.600 1082.240 ;
        RECT 4.400 1080.840 2695.600 1080.880 ;
        RECT 4.400 1079.480 2696.000 1080.840 ;
        RECT 3.990 1057.760 2696.000 1079.480 ;
        RECT 3.990 1056.400 2695.600 1057.760 ;
        RECT 4.400 1056.360 2695.600 1056.400 ;
        RECT 4.400 1055.000 2696.000 1056.360 ;
        RECT 3.990 1033.280 2696.000 1055.000 ;
        RECT 3.990 1031.920 2695.600 1033.280 ;
        RECT 4.400 1031.880 2695.600 1031.920 ;
        RECT 4.400 1030.520 2696.000 1031.880 ;
        RECT 3.990 1008.800 2696.000 1030.520 ;
        RECT 3.990 1007.440 2695.600 1008.800 ;
        RECT 4.400 1007.400 2695.600 1007.440 ;
        RECT 4.400 1006.040 2696.000 1007.400 ;
        RECT 3.990 985.680 2696.000 1006.040 ;
        RECT 3.990 984.280 2695.600 985.680 ;
        RECT 3.990 982.960 2696.000 984.280 ;
        RECT 4.400 981.560 2696.000 982.960 ;
        RECT 3.990 961.200 2696.000 981.560 ;
        RECT 3.990 959.800 2695.600 961.200 ;
        RECT 3.990 958.480 2696.000 959.800 ;
        RECT 4.400 957.080 2696.000 958.480 ;
        RECT 3.990 936.720 2696.000 957.080 ;
        RECT 3.990 935.320 2695.600 936.720 ;
        RECT 3.990 934.000 2696.000 935.320 ;
        RECT 4.400 932.600 2696.000 934.000 ;
        RECT 3.990 912.240 2696.000 932.600 ;
        RECT 3.990 910.840 2695.600 912.240 ;
        RECT 3.990 909.520 2696.000 910.840 ;
        RECT 4.400 908.120 2696.000 909.520 ;
        RECT 3.990 887.760 2696.000 908.120 ;
        RECT 3.990 886.360 2695.600 887.760 ;
        RECT 3.990 885.040 2696.000 886.360 ;
        RECT 4.400 883.640 2696.000 885.040 ;
        RECT 3.990 863.280 2696.000 883.640 ;
        RECT 3.990 861.880 2695.600 863.280 ;
        RECT 3.990 860.560 2696.000 861.880 ;
        RECT 4.400 859.160 2696.000 860.560 ;
        RECT 3.990 838.800 2696.000 859.160 ;
        RECT 3.990 837.400 2695.600 838.800 ;
        RECT 3.990 836.080 2696.000 837.400 ;
        RECT 4.400 834.680 2696.000 836.080 ;
        RECT 3.990 814.320 2696.000 834.680 ;
        RECT 3.990 812.920 2695.600 814.320 ;
        RECT 3.990 811.600 2696.000 812.920 ;
        RECT 4.400 810.200 2696.000 811.600 ;
        RECT 3.990 789.840 2696.000 810.200 ;
        RECT 3.990 788.440 2695.600 789.840 ;
        RECT 3.990 787.120 2696.000 788.440 ;
        RECT 4.400 785.720 2696.000 787.120 ;
        RECT 3.990 765.360 2696.000 785.720 ;
        RECT 3.990 763.960 2695.600 765.360 ;
        RECT 3.990 762.640 2696.000 763.960 ;
        RECT 4.400 761.240 2696.000 762.640 ;
        RECT 3.990 740.880 2696.000 761.240 ;
        RECT 3.990 739.480 2695.600 740.880 ;
        RECT 3.990 738.160 2696.000 739.480 ;
        RECT 4.400 736.760 2696.000 738.160 ;
        RECT 3.990 716.400 2696.000 736.760 ;
        RECT 3.990 715.000 2695.600 716.400 ;
        RECT 3.990 713.680 2696.000 715.000 ;
        RECT 4.400 712.280 2696.000 713.680 ;
        RECT 3.990 691.920 2696.000 712.280 ;
        RECT 3.990 690.520 2695.600 691.920 ;
        RECT 3.990 689.200 2696.000 690.520 ;
        RECT 4.400 687.800 2696.000 689.200 ;
        RECT 3.990 667.440 2696.000 687.800 ;
        RECT 3.990 666.040 2695.600 667.440 ;
        RECT 3.990 664.720 2696.000 666.040 ;
        RECT 4.400 663.320 2696.000 664.720 ;
        RECT 3.990 642.960 2696.000 663.320 ;
        RECT 3.990 641.560 2695.600 642.960 ;
        RECT 3.990 640.240 2696.000 641.560 ;
        RECT 4.400 638.840 2696.000 640.240 ;
        RECT 3.990 618.480 2696.000 638.840 ;
        RECT 3.990 617.080 2695.600 618.480 ;
        RECT 3.990 615.760 2696.000 617.080 ;
        RECT 4.400 614.360 2696.000 615.760 ;
        RECT 3.990 594.000 2696.000 614.360 ;
        RECT 3.990 592.600 2695.600 594.000 ;
        RECT 3.990 591.280 2696.000 592.600 ;
        RECT 4.400 589.880 2696.000 591.280 ;
        RECT 3.990 569.520 2696.000 589.880 ;
        RECT 3.990 568.120 2695.600 569.520 ;
        RECT 3.990 566.800 2696.000 568.120 ;
        RECT 4.400 565.400 2696.000 566.800 ;
        RECT 3.990 545.040 2696.000 565.400 ;
        RECT 3.990 543.640 2695.600 545.040 ;
        RECT 3.990 542.320 2696.000 543.640 ;
        RECT 4.400 540.920 2696.000 542.320 ;
        RECT 3.990 520.560 2696.000 540.920 ;
        RECT 3.990 519.160 2695.600 520.560 ;
        RECT 3.990 517.840 2696.000 519.160 ;
        RECT 4.400 516.440 2696.000 517.840 ;
        RECT 3.990 496.080 2696.000 516.440 ;
        RECT 3.990 494.680 2695.600 496.080 ;
        RECT 3.990 493.360 2696.000 494.680 ;
        RECT 4.400 491.960 2696.000 493.360 ;
        RECT 3.990 471.600 2696.000 491.960 ;
        RECT 3.990 470.200 2695.600 471.600 ;
        RECT 3.990 468.880 2696.000 470.200 ;
        RECT 4.400 467.480 2696.000 468.880 ;
        RECT 3.990 447.120 2696.000 467.480 ;
        RECT 3.990 445.720 2695.600 447.120 ;
        RECT 3.990 444.400 2696.000 445.720 ;
        RECT 4.400 443.000 2696.000 444.400 ;
        RECT 3.990 422.640 2696.000 443.000 ;
        RECT 3.990 421.240 2695.600 422.640 ;
        RECT 3.990 419.920 2696.000 421.240 ;
        RECT 4.400 418.520 2696.000 419.920 ;
        RECT 3.990 398.160 2696.000 418.520 ;
        RECT 3.990 396.760 2695.600 398.160 ;
        RECT 3.990 395.440 2696.000 396.760 ;
        RECT 4.400 394.040 2696.000 395.440 ;
        RECT 3.990 373.680 2696.000 394.040 ;
        RECT 3.990 372.280 2695.600 373.680 ;
        RECT 3.990 370.960 2696.000 372.280 ;
        RECT 4.400 369.560 2696.000 370.960 ;
        RECT 3.990 349.200 2696.000 369.560 ;
        RECT 3.990 347.800 2695.600 349.200 ;
        RECT 3.990 346.480 2696.000 347.800 ;
        RECT 4.400 345.080 2696.000 346.480 ;
        RECT 3.990 324.720 2696.000 345.080 ;
        RECT 3.990 323.320 2695.600 324.720 ;
        RECT 3.990 322.000 2696.000 323.320 ;
        RECT 4.400 320.600 2696.000 322.000 ;
        RECT 3.990 300.240 2696.000 320.600 ;
        RECT 3.990 298.840 2695.600 300.240 ;
        RECT 3.990 297.520 2696.000 298.840 ;
        RECT 4.400 296.120 2696.000 297.520 ;
        RECT 3.990 275.760 2696.000 296.120 ;
        RECT 3.990 274.360 2695.600 275.760 ;
        RECT 3.990 273.040 2696.000 274.360 ;
        RECT 4.400 271.640 2696.000 273.040 ;
        RECT 3.990 251.280 2696.000 271.640 ;
        RECT 3.990 249.880 2695.600 251.280 ;
        RECT 3.990 248.560 2696.000 249.880 ;
        RECT 4.400 247.160 2696.000 248.560 ;
        RECT 3.990 226.800 2696.000 247.160 ;
        RECT 3.990 225.400 2695.600 226.800 ;
        RECT 3.990 224.080 2696.000 225.400 ;
        RECT 4.400 222.680 2696.000 224.080 ;
        RECT 3.990 202.320 2696.000 222.680 ;
        RECT 3.990 200.920 2695.600 202.320 ;
        RECT 3.990 199.600 2696.000 200.920 ;
        RECT 4.400 198.200 2696.000 199.600 ;
        RECT 3.990 177.840 2696.000 198.200 ;
        RECT 3.990 176.440 2695.600 177.840 ;
        RECT 3.990 175.120 2696.000 176.440 ;
        RECT 4.400 173.720 2696.000 175.120 ;
        RECT 3.990 153.360 2696.000 173.720 ;
        RECT 3.990 151.960 2695.600 153.360 ;
        RECT 3.990 150.640 2696.000 151.960 ;
        RECT 4.400 149.240 2696.000 150.640 ;
        RECT 3.990 128.880 2696.000 149.240 ;
        RECT 3.990 127.480 2695.600 128.880 ;
        RECT 3.990 126.160 2696.000 127.480 ;
        RECT 4.400 124.760 2696.000 126.160 ;
        RECT 3.990 104.400 2696.000 124.760 ;
        RECT 3.990 103.000 2695.600 104.400 ;
        RECT 3.990 101.680 2696.000 103.000 ;
        RECT 4.400 100.280 2696.000 101.680 ;
        RECT 3.990 79.920 2696.000 100.280 ;
        RECT 3.990 78.520 2695.600 79.920 ;
        RECT 3.990 77.200 2696.000 78.520 ;
        RECT 4.400 75.800 2696.000 77.200 ;
        RECT 3.990 55.440 2696.000 75.800 ;
        RECT 3.990 54.040 2695.600 55.440 ;
        RECT 3.990 52.720 2696.000 54.040 ;
        RECT 4.400 51.320 2696.000 52.720 ;
        RECT 3.990 30.960 2696.000 51.320 ;
        RECT 3.990 29.560 2695.600 30.960 ;
        RECT 3.990 28.240 2696.000 29.560 ;
        RECT 4.400 26.840 2696.000 28.240 ;
        RECT 3.990 6.480 2696.000 26.840 ;
        RECT 3.990 5.080 2695.600 6.480 ;
        RECT 3.990 4.255 2696.000 5.080 ;
      LAYER met4 ;
        RECT 95.055 10.640 97.440 3457.360 ;
        RECT 99.840 10.640 2679.665 3457.360 ;
      LAYER met5 ;
        RECT 1168.060 2690.300 1170.580 2695.300 ;
  END
END ghazi_top_dffram_csv
END LIBRARY

